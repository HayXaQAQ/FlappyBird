// Verilog netlist created by TD v4.6.18154
// Sat Nov 14 16:17:28 2020

`timescale 1ns / 1ps
module moon  // al_ip/moon.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [13:0] addra;  // al_ip/moon.v(18)
  input clka;  // al_ip/moon.v(19)
  input rsta;  // al_ip/moon.v(20)
  output [7:0] doa;  // al_ip/moon.v(16)

  wire [0:1] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire \and_Naddra[12]_Naddr_o ;
  wire \and_Naddra[12]_addra_o ;
  wire \and_addra[12]_Naddra_o ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  and \and_Naddra[12]_Naddr  (\and_Naddra[12]_Naddr_o , ~addra[12], ~addra[13]);
  and \and_Naddra[12]_addra  (\and_Naddra[12]_addra_o , ~addra[12], addra[13]);
  and \and_addra[12]_Naddra  (\and_addra[12]_Naddra_o , addra[12], ~addra[13]);
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_01(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_02(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_03(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_04(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_05(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_06(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_07(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_08(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_09(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0A(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0C(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0D(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0F(256'h808080808080808080808080808080808080808080808080808080808080B3B3),
    .INIT_10(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_11(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_12(256'h8080808080808080808080808080808080808080808080808080B3B380808080),
    .INIT_13(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_14(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_15(256'h808080808080808080808080808080808080808080B3B3B38080808080808080),
    .INIT_16(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_17(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_18(256'h80808080808080808080808080808080B3B3B3B3808080808080808080808080),
    .INIT_19(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1A(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1B(256'h8080808080808080808080B3B3B3B3B380808080808080808080808080808080),
    .INIT_1C(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1D(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1E(256'h808080808080B3B3B3B3B3B3B380808080808080808080808080808080808080),
    .INIT_1F(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_20(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_21(256'h8080B3B3B3B3B3B3B38080808080808080808080808080808080808080808080),
    .INIT_22(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_23(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_24(256'hB3B3B3B3B3808080808080808080808080808080808080808080808080808080),
    .INIT_25(256'h8080808080808080808080808080808080808080808080808080808080B3B3B3),
    .INIT_26(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_27(256'hB380808080808080808080808080808080808080808080808080808080808080),
    .INIT_28(256'h808080808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3),
    .INIT_29(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_2A(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_2B(256'h8080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3808080),
    .INIT_2C(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_2D(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_2E(256'h808080808080808080808080808080B3B3B3B3B3B3B3B3B3B380808080808080),
    .INIT_2F(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_30(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_31(256'h8080808080808080808080B3B3B3B3B3B3B3B3B3B38080808080808080808080),
    .INIT_32(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_33(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_34(256'h808080808080B3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080),
    .INIT_35(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_36(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_37(256'h8080B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080808080),
    .INIT_38(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_39(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_3A(256'hB3B3B3B3B3B3B3B3B3B380808080808080808080808080808080808080808080),
    .INIT_3B(256'h8080808080808080808080808080808080808080808080808080808080B3B3B3),
    .INIT_3C(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_3D(256'hB3B3B3B3B3B38080808080808080808080808080808080808080808080808080),
    .INIT_3E(256'h80808080808080808080808080808080808080808080808080B3B3B3B3B3B3B3),
    .INIT_3F(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_40(256'hB3B3808080808080808080808080808080808080808080808080808080808080),
    .INIT_41(256'h8080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_42(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_43(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_44(256'h80808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B38080),
    .INIT_45(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_46(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_47(256'h8080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080),
    .INIT_48(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_49(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_4A(256'h80808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080),
    .INIT_4B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_4C(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_4D(256'h808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080808080808080808080),
    .INIT_4E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_4F(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_50(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080808080),
    .INIT_51(256'h808080808080808080808080808080808080808080808080808080808080B3B3),
    .INIT_52(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_53(256'hB3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080808080808080),
    .INIT_54(256'h8080808080808080808080808080808080808080808080808080B3B3B3B3B3B3),
    .INIT_55(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_56(256'hB3B3B3B3B3B3B3B3808080808080808080808080808080808080808080808080),
    .INIT_57(256'h80808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3),
    .INIT_58(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_59(256'hB3B3B3B380808080808080808080808080808080808080808080808080808080),
    .INIT_5A(256'h8080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_5B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_5C(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_5D(256'h80808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_5E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_5F(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_60(256'h808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080),
    .INIT_61(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_62(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_63(256'h8080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080808080),
    .INIT_64(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_65(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_66(256'h80B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080),
    .INIT_67(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_68(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_69(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080),
    .INIT_6A(256'h80808080808080808080808080808080808080808080808080808080B3B3B3B3),
    .INIT_6B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_6C(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080808080),
    .INIT_6D(256'h808080808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3),
    .INIT_6E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_6F(256'hB3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080808080808080),
    .INIT_70(256'h8080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_71(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_72(256'hB3B3B3B3B3B3B380808080808080808080808080808080808080808080808080),
    .INIT_73(256'h80808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_74(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_75(256'hB3B3B3B380808080808080808080808080808080808080808080808080808080),
    .INIT_76(256'h808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_77(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_78(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_79(256'h80808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_7A(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_7B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_7C(256'h808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080),
    .INIT_7D(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_7E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_7F(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080808080),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_10000x8_sub_000000_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_Naddra[12]_Naddr_o ),
    .dia({open_n51,open_n52,open_n53,open_n54,open_n55,open_n56,open_n57,open_n58,8'b00000000}),
    .rsta(rsta),
    .doa({open_n80,open_n81,open_n82,open_n83,open_n84,open_n85,open_n86,open_n87,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=4096;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h80808080808080808080808080808080808080808080808080808080808080B3),
    .INIT_01(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_02(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080808080808080),
    .INIT_03(256'h808080808080808080808080808080808080808080808080808080B3B3B3B3B3),
    .INIT_04(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_05(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080),
    .INIT_06(256'h8080808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3),
    .INIT_07(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_08(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080808080),
    .INIT_09(256'h80808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_0A(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0B(256'hB3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080808080808080),
    .INIT_0C(256'h808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_0D(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0E(256'hB3B3B3B3B3B3B3B3808080808080808080808080808080808080808080808080),
    .INIT_0F(256'h8080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_10(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_11(256'hB3B3B3B380808080808080808080808080808080808080808080808080808080),
    .INIT_12(256'h8080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_13(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_14(256'hB380808080808080808080808080808080808080808080808080808080808080),
    .INIT_15(256'h80808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_16(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_17(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_18(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080),
    .INIT_19(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1A(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1B(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080),
    .INIT_1C(256'h80808080808080808080808080808080808080808080808080808080B3B3B3B3),
    .INIT_1D(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1E(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080),
    .INIT_1F(256'h808080808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3),
    .INIT_20(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_21(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080808080),
    .INIT_22(256'h8080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_23(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_24(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080),
    .INIT_25(256'h80808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_26(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_27(256'hB3B3B3B3B3B3B3B3B3B3B3B3B380808080808080808080808080808080808080),
    .INIT_28(256'h80808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_29(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_2A(256'hB3B3B3B3B3B3B3B3B3B380808080808080808080808080808080808080808080),
    .INIT_2B(256'h808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_2C(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_2D(256'hB3B3B3B3B3B3B380808080808080808080808080808080808080808080808080),
    .INIT_2E(256'h8080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_2F(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_30(256'hB3B3B3B380808080808080808080808080808080808080808080808080808080),
    .INIT_31(256'h80B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_32(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_33(256'hB380808080808080808080808080808080808080808080808080808080808080),
    .INIT_34(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_35(256'h808080808080808080808080808080808080808080808080808080808080B3B3),
    .INIT_36(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_37(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080),
    .INIT_38(256'h8080808080808080808080808080808080808080808080808080B3B3B3B3B3B3),
    .INIT_39(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_3A(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080),
    .INIT_3B(256'h80808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3),
    .INIT_3C(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_3D(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080),
    .INIT_3E(256'h80808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_3F(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_40(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080),
    .INIT_41(256'h808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_42(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_43(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080),
    .INIT_44(256'h808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_45(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_46(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080808080),
    .INIT_47(256'h8080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_48(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_49(256'hB3B3B3B3B3B3B3B3B3B3B3B3B380808080808080808080808080808080808080),
    .INIT_4A(256'h80808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_4B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_4C(256'hB3B3B3B3B3B3B3B3B3B380808080808080808080808080808080808080808080),
    .INIT_4D(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_4E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_4F(256'hB3B3B3B3B3B3B380808080808080808080808080808080808080808080808080),
    .INIT_50(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_51(256'h8080808080808080808080808080808080808080808080808080808080B3B3B3),
    .INIT_52(256'hB3B3B3B380808080808080808080808080808080808080808080808080808080),
    .INIT_53(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_54(256'h8080808080808080808080808080808080808080808080808080B3B3B3B3B3B3),
    .INIT_55(256'hB380808080808080808080808080808080808080808080808080808080808080),
    .INIT_56(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_57(256'h80808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3),
    .INIT_58(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_59(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380),
    .INIT_5A(256'h80808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_5B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_5C(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080),
    .INIT_5D(256'h808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_5E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_5F(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080),
    .INIT_60(256'h808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_61(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_62(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080),
    .INIT_63(256'h8080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_64(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_65(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080),
    .INIT_66(256'h8080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_67(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_68(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080),
    .INIT_69(256'h8080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_6A(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_6B(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080808080808080808080),
    .INIT_6C(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_6D(256'h808080808080808080808080808080808080808080808080808080808080B3B3),
    .INIT_6E(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080),
    .INIT_6F(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_70(256'h808080808080808080808080808080808080808080808080808080B3B3B3B3B3),
    .INIT_71(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080808080808080808080808080),
    .INIT_72(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_73(256'h808080808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3),
    .INIT_74(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080808080),
    .INIT_75(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_76(256'h808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_77(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080808080),
    .INIT_78(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_79(256'h8080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_7A(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080808080),
    .INIT_7B(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_7C(256'h808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_7D(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080808080808080808080808080),
    .INIT_7E(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_7F(256'h808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_10000x8_sub_004096_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_addra[12]_Naddra_o ),
    .dia({open_n108,open_n109,open_n110,open_n111,open_n112,open_n113,open_n114,open_n115,8'b00000000}),
    .rsta(rsta),
    .doa({open_n137,open_n138,open_n139,open_n140,open_n141,open_n142,open_n143,open_n144,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  // address_offset=8192;data_offset=0;depth=1808;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080),
    .INIT_01(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_02(256'h8080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_03(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080808080808080),
    .INIT_04(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_05(256'h8080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_06(256'hB3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080808080808080),
    .INIT_07(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_08(256'h8080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_09(256'hB3B3B3B3B3B3B380808080808080808080808080808080808080808080808080),
    .INIT_0A(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_0B(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_0C(256'hB3B38080808080808080808080808080808080808080808080808080808080B3),
    .INIT_0D(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_0E(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_0F(256'h8080808080808080808080808080808080808080808080808080808080B3B3B3),
    .INIT_10(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080),
    .INIT_11(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_12(256'h8080808080808080808080808080808080808080808080808080B3B3B3B3B3B3),
    .INIT_13(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3808080808080808080),
    .INIT_14(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_15(256'h808080808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3),
    .INIT_16(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080),
    .INIT_17(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_18(256'h808080808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_19(256'hB3B3B3B3B3B3B3B3B3B3B3B38080808080808080808080808080808080808080),
    .INIT_1A(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_1B(256'h80808080808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_1C(256'hB3B3B3B3B3B38080808080808080808080808080808080808080808080808080),
    .INIT_1D(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_1E(256'h80808080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_1F(256'hB380808080808080808080808080808080808080808080808080808080808080),
    .INIT_20(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_21(256'h8080808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_22(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_23(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080808080),
    .INIT_24(256'h808080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_25(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_26(256'hB3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B380808080808080808080808080),
    .INIT_27(256'h8080808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_28(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_29(256'hB3B3B3B3B3B3B3B3B3B3B3B3B380808080808080808080808080808080808080),
    .INIT_2A(256'h808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_2B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_2C(256'hB3B3B3B3B3B38080808080808080808080808080808080808080808080808080),
    .INIT_2D(256'h8080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_2E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_2F(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_30(256'h808080808080808080B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B38080),
    .INIT_31(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_32(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_33(256'h8080808080808080808080B3B3B3B3B3B3B3B3B3808080808080808080808080),
    .INIT_34(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_35(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_36(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_37(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_38(256'h0000000000000000000000000000000080808080808080808080808080808080),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_10000x8_sub_008192_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(\and_Naddra[12]_addra_o ),
    .dia({open_n165,open_n166,open_n167,open_n168,open_n169,open_n170,open_n171,open_n172,8'b00000000}),
    .rsta(rsta),
    .doa({open_n194,open_n195,open_n196,open_n197,open_n198,open_n199,open_n200,open_n201,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i2_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i2_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i2_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i2_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i2_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i2_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i2_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i2_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[7]));

endmodule 

