// Verilog netlist created by TD v4.6.18154
// Wed Nov 11 23:53:02 2020

`timescale 1ns / 1ps
module Startbutton  // al_ip/Startbutton.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [12:0] addra;  // al_ip/Startbutton.v(18)
  input clka;  // al_ip/Startbutton.v(19)
  input rsta;  // al_ip/Startbutton.v(20)
  output [7:0] doa;  // al_ip/Startbutton.v(16)

  wire [0:0] addra_piped;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;

  reg_sr_as_w1 addra_pipe (
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSAMUX("INV"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'hA7A7A7A7A7A7A7A7A7A7A7A7A7A7A7A8A8A8A7A6A6A6A7A7A5A7A3A4A39D908B),
    .INIT_01(256'hA8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A7A7A7A7A7A7A7A7A7A7A7A7A7A7A7A7A7),
    .INIT_02(256'hA8A8A7A7A8A8A8A7A8A8A8A8A8A8A7A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8),
    .INIT_03(256'h8E8E8E8E8E8E8E8E8E8E8E8E8E8F8F8F8E8E90908E908A8F90928989B9AAA4A5),
    .INIT_04(256'h91919191919191919191919191909090909090908E8E8E8E8E8E8E8E8E8E8E8E),
    .INIT_05(256'h909090919191929191908F909091919191919191919191919191919191919191),
    .INIT_06(256'h8D8D8D8D8D8D8D8C8C8C8D8D8C8C8E8E8B8B868A8A8E8B8CAA958E919292908F),
    .INIT_07(256'h8C8C8C8C8C8C8C8C8B8C8C8B8B8B8B8B8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D),
    .INIT_08(256'h8C8D8D8D8C8C8A8B8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C),
    .INIT_09(256'h91919191909091918F909292939491938D8D8A8AA88F888A8D8C8B8C8B8B8B8C),
    .INIT_0A(256'h9292929293939392929292929191919191919191919191919191919191919191),
    .INIT_0B(256'h9292919192929292929292929292929292929292929292929292929292929292),
    .INIT_0C(256'h9C9C9B9B9B9B9D9D9A9B9B9A8F8E8989A8918B8E919192929292919292929292),
    .INIT_0D(256'h999999999A9A9A9A9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9C),
    .INIT_0E(256'h9898979897989798979897989798979897989798979897989798979897989798),
    .INIT_0F(256'h9E9FA1A1A2A1A19F8E8C8A8AA58E8C9094969897979897979798989898979797),
    .INIT_10(256'hA0A1A1A19F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9FA0A0A09E9E),
    .INIT_11(256'h9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9FA0A0A0),
    .INIT_12(256'hA2A1A19E8A878787A48F8C919A9D9F9F9E9E9F9E9E9F9F9F9E9E9E9E9E9F9F9F),
    .INIT_13(256'hA1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A0A0A0A1A2A2),
    .INIT_14(256'hA1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A0A0A0A0A0A0A0A0),
    .INIT_15(256'h8B898B8BA38D8C929B9FA3A2A0A1A2A0A1A2A2A2A1A1A1A1A1A1A1A1A1A1A1A1),
    .INIT_16(256'hA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A09F9F9E9FA0A09F9FA09E),
    .INIT_17(256'hA1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A0A0A0A0A0A0A0A0A0),
    .INIT_18(256'hA48F8E939A9EA2A1A0A0A09FA1A1A1A1A1A1A0A0A1A1A1A1A1A1A1A1A1A1A1A1),
    .INIT_19(256'hA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A09F9F9F9FA0A09F9F9F9D8E8A898A),
    .INIT_1A(256'hA1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0),
    .INIT_1B(256'h9B9FA2A1A1A19FA0A1A1A1A1A1A1A0A0A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1),
    .INIT_1C(256'hA0A0A0A0A0A0A0A0A0A0A0A0A1A1A0A09F9FA1A09F9F9F9D8E8B8A8AA48D8B92),
    .INIT_1D(256'hA1A0A1A0A1A0A1A0A1A0A1A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0),
    .INIT_1E(256'hA0A09FA0A1A0A0A0A0A1A0A0A1A0A1A0A1A0A1A0A1A0A1A0A1A0A1A0A1A0A1A0),
    .INIT_1F(256'hA1A1A1A1A1A1A1A1A1A2A2A1A09FA0A19FA0A09E8D8A8A8CA48D8B929A9FA2A1),
    .INIT_20(256'hA0A0A0A0A0A0A0A0A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1),
    .INIT_21(256'hA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0),
    .INIT_22(256'hA1A1A1A1A1A1A2A2A0A0A1A19FA1A09E8D8A8A8CA48D8B919A9FA2A0A0A09FA0),
    .INIT_23(256'hA0A0A0A0A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1),
    .INIT_24(256'hA0A09F9FA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0),
    .INIT_25(256'hA1A1A1A2A1A1A1A1A0A09F9E8D8A8A8CA48D8B919A9EA2A0A0A09E9F9FA0A0A0),
    .INIT_26(256'hA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A1),
    .INIT_27(256'hA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0),
    .INIT_28(256'hA1A1A2A19F9F9F9D8C8A8A8CA48D8B91999EA19F9F9F9E9F9F9F9F9F9F9F9F9F),
    .INIT_29(256'hA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A1),
    .INIT_2A(256'hA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0),
    .INIT_2B(256'h9F9F9E9C8D898A8CA48C8A91999EA1A0A09F9E9F9FA09FA09F9FA0A0A0A0A0A0),
    .INIT_2C(256'hA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A09F9F9F9F9FA0A0A1A1),
    .INIT_2D(256'hA0A1A0A1A0A1A0A1A0A1A0A1A0A1A0A1A0A1A0A1A0A1A0A0A0A0A0A0A0A0A0A0),
    .INIT_2E(256'h8C898A8CA38C8A919A9FA2A1A1A09FA0A0A0A0A1A0A0A0A0A0A1A0A1A0A1A0A1),
    .INIT_2F(256'hA7A7A7A7A6A6A6A5A4A4A4A4A4A5A5A6A7A7A7A7A6A5A3A3A1A1A1A09FA09F9D),
    .INIT_30(256'hA9AAAAA9A9A8A8A7A6A4A2A0A0A0A1A2A3A5A8A7A6A4A1A0A1A2A3A5A6A7A7A8),
    .INIT_31(256'hA38C8A919AA0A4A4A6A7A7A8A8A8A7A7A7A7A6A6A6A6A5A5A5A5A3A3A4A5A6A8),
    .INIT_32(256'hA7A8ABAAABAAA6A9A8B1ABA6A9A5A4A7A7A6A7A7A6A2A0A0A1A2A09D8D8A8B8C),
    .INIT_33(256'hA9ABA8A9A3A8A3A09FA19F9FA8AEABA4A6A7A5A29FA9ADA9A6A6A3A8A7A7ACA8),
    .INIT_34(256'h98A0A5ACAEA7A4A3A6A5A6A6A7ACADA8ACABABAAAAA8A6A7A9ABABA8A7A8A8A8),
    .INIT_35(256'hA1A09A9FA4B2ADA2A6A7A6A3A3A3A2A5A6A5A3A0A1A2A19D8D8A8B8CA38D8B91),
    .INIT_36(256'h9FA7A29F9DA1A1A5B1B5B1A7A5A6A5A4A2A8AEAFA2A5A4A9A8A7A9A1A6A4A5A3),
    .INIT_37(256'hADA4A3A2A4A5A7A6A4A5A7A3A3A1A19F9EA2A8AEB0AAA1A0A6A8A7A7AAAAA5A5),
    .INIT_38(256'hAFBCB2A2A7B1B6B5B3AFA59FA1A6A3A19FA1A09D8C898A8CA48D8B919AA1A6AB),
    .INIT_39(256'h9EA1A2ABBABEB3A7A4A4A7A9A7A7AFB1ABAFB0B4B8BAB8ACA8A6A9A9A7A59EA2),
    .INIT_3A(256'hB2B5B9BAB3AAA8AAA7A7A8A29BA1ADB8B9ADA2A8B1B2B3B8B6B4A7A19DA8A29E),
    .INIT_3B(256'hA9B4BABCC2C2B8A8A1A4A3A29F9FA09D8B888A8CA38D8B929EA5A9AFB2AEB0B0),
    .INIT_3C(256'hC0C1B3A9ACA6A6ABA8A7ACAEAEB2B2B8BFC4C6BBADADB6BBB9B5AFB0B6BEB4A5),
    .INIT_3D(256'hC1B1ACB2B6B7B8B1A8ABB7C0B7ABA6B2B6B5B5BFC5C3B2A6A0ABA49EA0A2A3AF),
    .INIT_3E(256'hBAC3C2B8ABA7A5A5A1A0A09D8A878A8DA38D8B929BA3A7ADB1AFB1B3B6BAC2C5),
    .INIT_3F(256'hB4A9A3A6A6A4A5A6A3A8A7ACB5BFC6BCAEAAB2B7B5B2ADAFB1B6B0ABA9AAAEAD),
    .INIT_40(256'hB4B2B2B0ACB1BCC4B8A9A4ADAEAAAAB4C6C7B5A7A1ACA5A0A1A4A9B5C3BCAFAB),
    .INIT_41(256'hACA5A3A6A1A0A19D8A878A8DA38D8B919BA2A3A5A7A3A5A6A9B0BCC5C2B0AAB1),
    .INIT_42(256'hA6A5A2A2A0A3A1A6AFBBC7C2B1A6ACAFABA9A6A7ACACAAA9A7A7ACAEB8C2C4B9),
    .INIT_43(256'hA6AEBAC2BEB0A5A9ABABA9B1C3C8B9AAA1ACA6A0A1A6AFBCC3B6AAADBCB4A6A2),
    .INIT_44(256'hA2A3A39F8C898B8DA38D8B919BA1A2A3A3A0A0A0A2ABB8C3C4B3A8ACAEA9A9A7),
    .INIT_45(256'hA0A3A2A7ADB8C7C7B6A6A7ABA4A2A1A2A1A29FA3A2A4ACB0B8BEBBB2A7A2A2A5),
    .INIT_46(256'hBFB7ABA7A9ACACB3C1C7BCAEA0ACA7A2A2A8B4BEBEAEA7B1C3C0B1A4A8ABA4A2),
    .INIT_47(256'h8D898A8CA38D8B90959D9EA0A2A09F9EA0A9B5C0C5B4A4A4A9A4A4A2A1A9B5BC),
    .INIT_48(256'hABB4C4C6B5A4A6A9A19E9D9FA0A6A6AAA8A9AFACAEAFACA9A5A4A2A5A2A3A39F),
    .INIT_49(256'hA3A8AEB4BEC4BCADA0AAA7A3A3ABB8C0BBA9AAB8C6C6BAA6AAAEA6A29FA0A0A6),
    .INIT_4A(256'hA38D8B91999FA1A3A3A09F9C9FA8B1BEC6B8A7A3A7A2A3A1A1A7B0B6C0BFB7A9),
    .INIT_4B(256'hB6A7A2A8A09A9B9FA4A9ACAEAEACA9A7ABA5A7A8A3A5A5A2A2A3A29E8C89898B),
    .INIT_4C(256'hAEB8BCB4A4A6A5A4A6B0BFC3B6ABB1BBC8C5BCAFA8A9A8A6A09E9EA2A7B3C0C7),
    .INIT_4D(256'h9A9FA2A1A3A29F9FA1A6B3BDC8BAADA3A6A4A1A1A4A2A7AFB6BCBEBCB2AAA8AD),
    .INIT_4E(256'hA19B9DA2A8B0B3B0ABA9AAA9AAA7ADAFA9A5A29CA2A3A19D8C88888AA38D8B91),
    .INIT_4F(256'hA6A8A6A6A7B5C1BFB2ACAFB3B7BAB9B3ACA9A9A9A39F9E9FA4AFBFC8B4A5A1A9),
    .INIT_50(256'hA3A3A0A0A0A3B1BBC7BAAEA3A7A5A3A2A5A1A2A8B0B7BFC2BFB7ADA8A9B4BBB2),
    .INIT_51(256'hB2BABAAFA6A7ABABADAAABA9A5A4A39EA4A5A19C8B88888AA38D8B919B9FA2A1),
    .INIT_52(256'hAEBCC1B7ADB0B0ADADADAEAEADACA8A4A9A4A09FA2AEC1CBB6A6A3ABA5A0A3A8),
    .INIT_53(256'h9EA3AFBBC7BBB0A6A7A4A1A0A2A0A2A5AEB5BBBEBDB5AAA6B3BAC0B4A8A8A7A8),
    .INIT_54(256'hA8AFB2B1AFAAA69F9C9EA1A1A4A5A19D8C89898AA38D8B919B9EA09FA1A2A0A0),
    .INIT_55(256'hAAB4B5B2B5B1ACAEB0ADA9A2ABA6A4A2A1ABC1CDB8A7A4ADA7A3A5AAB8BFBCAE),
    .INIT_56(256'hC8BCB1A7A8A39F9EA0A3A6AAB1B5B5B0ACA8A9AEBBC1C5B6A9A6A9ADB8C0BDAE),
    .INIT_57(256'hADAAA6A3A2A2A2A2A4A5A29F8E8B8B8CA38D8B929B9FA09EA0A0A0A09EA3AFBB),
    .INIT_58(256'hB4B8BAB9B7B0ACA6A8A7A6A4A3ABC0CDB8A6A1ABA6A0A2A8B7BFBFB3AAACB0B0),
    .INIT_59(256'hA9A4A0A0A2A7AEAEB2B1ACA6A5A6A7AEB6BFC5B4A8A5AEB3BDBDB2A7A7B1B3B3),
    .INIT_5A(256'hA7A5A4A7A4A3A19E8E8B8B8DA38D8B929CA0A09EA0A0A0A0A0A3B1BCC8BBAFA5),
    .INIT_5B(256'hC0BDB3A5A2A4A5A3A3ABC0CCB6A59FA9A5A0A1A5B0BDC2BCADA5A6A7A7A8A5A5),
    .INIT_5C(256'hA6ACB3ADA8A5A3A5ABABA5A7B0BDC7B4AAA6B3B9BEB5A9A4A6ACADAFAFB4B8BD),
    .INIT_5D(256'hA4A19F9B8C8A8B8DA38D8B929DA1A09D9FA0A0A0A1A4B0BBC7B8AAA1A6A2A2A3),
    .INIT_5E(256'hA2A5A5A3A4ACC0C9B6A5A0A9A6A1A0A3A9B5BDBDB6AEACAEA9A7A4A5A8A49FA7),
    .INIT_5F(256'hA8A7A7ABAAA6A1A2B1BFCAB6ACA8B9BEBAB0A9AAA9A8A4A4A5A8ABB4C2C6BBA8),
    .INIT_60(256'h8B898A8CA38D8B929DA09F9D9E9F9FA0A1A3B0BBC6B8AAA1A4A1A4A8ABB3BCB0),
    .INIT_61(256'hA4ABBAC2B1A29FA8A6A1A0A1A8ABB2B9BBB8B7B5ADACA6A8A89D9AA6A5A19E9A),
    .INIT_62(256'hA6A09EA3B2BDC5ACA5A4BAC1AFA9A6A9ABA8A19C9CA2A7ABB9C0BBAF9FA3A4A3),
    .INIT_63(256'hA38D8B929B9FA09D9FA09FA1A0A2ADB6C0B2A49FA3A1A5A9ABB5BCAEA7AAADAC),
    .INIT_64(256'hAEABA8A4A2A1A0A2A1A6ACB0B4B7B9BBB6B2ADA7A39FA3A5A5A29F9B8A88888A),
    .INIT_65(256'hAEB9B8ADA2A6B3BAAFA9A7A8A7A3A0A09FA2A5AAAFB2B2B0A7A4A2A3A6AAB0B3),
    .INIT_66(256'h9CA0A1A0A0A1A0A2A2A5A9ACADADAAA5A4A1A3A6A9ACB0B2ACACAAA7A5A1A0A4),
    .INIT_67(256'hA0A09F9FA0A2A6A9ACAEB0B3B5B4B2AFABA7A6A7A4A2A09D8B88898BA38D8B91),
    .INIT_68(256'hA7AAB0B1ADA7A4A5A5A2A0A09EA0A3A6A8A9A9A7A1A1A0A2A4A6A7A8A6A5A5A3),
    .INIT_69(256'hA1A0A0A2A1A3A4A6A6A5A5A2A1A0A2A4A6A7A8A8A4A4A3A3A1A09EA2AAB2B2AD),
    .INIT_6A(256'h9FA0A1A3A5A6A8AAABAAAAACA9A5A4A4A1A1A09E8E8C8D8EA38E8B909B9FA1A0),
    .INIT_6B(256'hA8A5A4A4A3A09E9F9D9D9FA1A3A4A3A2A1A09FA0A0A2A3A3A4A2A2A09F9F9E9E),
    .INIT_6C(256'hA0A2A2A3A4A4A4A29F9FA0A1A2A3A4A4A3A2A2A19F9E9D9EA0A6A8A7A7A8A8A6),
    .INIT_6D(256'hA0A0A2A3A3A1A1A2A2A1A1A1A0A1A09E8E8D8D8EA38E8B909B9FA1A09FA09FA1),
    .INIT_6E(256'hA09E9E9F9D9D9E9FA0A0A0A0A09F9F9F9FA0A1A1A0A0A0A09FA0A0A0A09FA0A0),
    .INIT_6F(256'hA1A1A1A19F9FA0A0A2A2A2A2A1A0A09F9F9F9F9F9C9E9F9FA1A3A29FA2A1A1A2),
    .INIT_70(256'hA09E9EA0A1A1A2A2A0A1A09D8E8B8B8CA38E8B909B9FA1A09F9F9EA1A1A1A2A1),
    .INIT_71(256'h9F9F9F9F9FA0A0A1A1A0A0A0A1A0A1A19F9FA0A1A1A2A2A2A1A1A0A09F9E9E9E),
    .INIT_72(256'hA1A1A2A2A2A2A2A1A19F9F9FA1A1A2A19F9F9E9D9EA0A09F9F9FA0A0A09FA0A1),
    .INIT_73(256'hA1A2A2A2A0A1A09D8D8A898AA38E8B919BA0A2A1A0A09EA0A1A1A0A09F9F9FA0),
    .INIT_74(256'h9F9FA0A1A2A2A2A2A0A09F9F9FA0A0A1A1A2A2A2A1A2A1A09F9E9C9C9D9EA0A0),
    .INIT_75(256'hA2A1A1A0A0A0A0A0A0A2A2A2A1A0A19F9F9F9F9F9E9E9E9F9F9F9FA0A1A1A0A0),
    .INIT_76(256'hA0A1A09D8C898889A38E8B919CA1A2A2A0A09FA19FA0A09FA0A09FA0A1A2A2A2),
    .INIT_77(256'hA2A2A3A2A2A09F9F9FA0A0A0A1A1A1A1A1A1A1A0A0A0A09F9D9FA0A0A0A1A1A0),
    .INIT_78(256'h9F9F9FA0A0A1A2A2A2A2A2A2A0A09F9F9E9E9E9E9E9E9E9FA2A2A1A09F9FA0A1),
    .INIT_79(256'h8D89898AA38E8B919CA1A3A2A1A09FA1A0A0A0A0A0A09FA0A0A1A1A1A0A0A09F),
    .INIT_7A(256'hA2A1A09F9F9FA0A0A0A1A1A1A0A0A1A0A1A1A2A2A0A1A1A1A0A0A2A2A0A1A09D),
    .INIT_7B(256'hA1A1A1A2A3A2A2A2A1A0A0A1A0A09F9FA0A1A0A0A2A2A1A09F9FA0A0A2A2A3A3),
    .INIT_7C(256'hA38E8B919CA1A3A2A1A09FA1A1A1A1A1A1A0A09FA0A0A0A0A0A09F9F9F9F9FA0),
    .INIT_7D(256'hA0A0A0A0A0A09FA0A0A0A1A1A2A2A2A2A1A1A1A1A1A1A1A19F9FA29D908B8C8B),
    .INIT_7E(256'hA1A1A1A1A1A1A2A2A2A2A1A1A1A2A2A2A1A1A1A1A0A0A0A1A1A2A2A1A1A0A0A0),
    .INIT_7F(256'h9DA1A29F9F9F9FA0A1A1A1A1A1A0A0A09F9F9FA0A0A0A0A0A09F9F9FA0A0A0A1),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_5000x8_sub_000000_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(addra[12]),
    .dia({open_n51,open_n52,open_n53,open_n54,open_n55,open_n56,open_n57,open_n58,8'b00000000}),
    .rsta(rsta),
    .doa({open_n80,open_n81,open_n82,open_n83,open_n84,open_n85,open_n86,open_n87,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=4096;data_offset=0;depth=904;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h9F9F9F9F9FA0A0A0A1A2A2A2A2A1A1A19F9FA0A09E9FA29D908A8D8DA48E898E),
    .INIT_01(256'hA0A1A1A2A2A2A2A2A2A2A1A1A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0),
    .INIT_02(256'h9F9F9EA0A0A0A0A0A0A0A09F9F9E9FA0A0A0A0A0A0A0A09F9F9FA09F9F9F9FA0),
    .INIT_03(256'hA0A0A0A0A0A0A0A1A1A1A1A19F9FA1A1A09FA29D908A8C8CA48E898E9CA0A19E),
    .INIT_04(256'hA1A2A2A2A1A1A1A0A0A0A0A1A1A1A1A1A0A09F9FA0A0A0A1A1A1A1A1A1A1A1A0),
    .INIT_05(256'hA0A0A1A1A1A1A1A09F9FA0A1A2A3A3A3A2A2A1A1A0A0A0A09E9E9E9FA0A0A1A2),
    .INIT_06(256'hA1A0A1A1A3A3A3A2A0A1A1A1A0A0A19D918A8C8AA48E8A8E9DA0A19FA09F9EA0),
    .INIT_07(256'hA2A1A1A1A0A1A1A2A2A2A2A2A1A0A1A0A1A1A2A2A2A2A2A2A2A2A2A2A2A2A1A1),
    .INIT_08(256'hA3A2A2A2A1A1A2A2A4A4A4A4A4A3A3A2A2A2A2A19F9E9FA0A0A1A2A2A2A3A2A2),
    .INIT_09(256'h9FA09F9E9E9E9F9F9F9EA09B908B8B89A48F8A8D9EA1A2A1A1A1A0A1A2A2A2A2),
    .INIT_0A(256'h9E9FA0A0A1A0A0A0A09F9F9FA0A0A1A0A1A0A1A0A1A1A1A1A1A0A0A09F9E9E9E),
    .INIT_0B(256'hA0A0A1A1A2A2A2A2A2A1A1A0A1A0A1A09E9E9E9E9E9F9F9F9F9F9E9E9E9E9E9E),
    .INIT_0C(256'h98999A9A9A989A978E8B8B87A38F8A8C9EA1A1A0A1A09FA1A2A2A2A2A2A2A2A1),
    .INIT_0D(256'h9B9B9B9A9A9A9A9A9B9B9B9B9B9B9B9B9B9B9B9B9B9B9A9A9999999999999998),
    .INIT_0E(256'h9B9B9B9B9B9A9A9A9B9B9B9B9A9A9A99999999999999999898989999999A9A9B),
    .INIT_0F(256'h938F91928C8B8C89A38F898B999C9B9B9B9A999B9C9C9C9C9C9C9B9B9B9B9B9B),
    .INIT_10(256'h9393939394949493939292929292929292929393939394939292929291939393),
    .INIT_11(256'h9191919192939394939394939392919191919192939393939393939393939393),
    .INIT_12(256'h8A8C8D89A490888B9193929192918F9292929292929190919293939393929291),
    .INIT_13(256'h8B8B8B8A8A8A8A898989898989898A8A8B8B8C8B8A8A8A8A8A8A8C8B8B878A8D),
    .INIT_14(256'h898A8A8B8B8B8B8B8A8A898989898A8A8B8B8C8B8B8B8A8A8A8A8A8A8A8B8B8B),
    .INIT_15(256'hA490898A8A8C8B898B89888B89898989888888888A8A8A8A8A89898888888888),
    .INIT_16(256'h8B8B8B8A8A8A8A8A8A8A8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8A8A8B8C8C8C8B),
    .INIT_17(256'h8B8B8B8B8B8B8A8A8A8A8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B),
    .INIT_18(256'h8B8B8B8A8A8A8A8A8A8A8A8A8A8A8A8A8B8B8B8B8B8A8A8A8A8A8A8A8A8B8B8B),
    .INIT_19(256'h8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8CA38F8B8B),
    .INIT_1A(256'h8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C),
    .INIT_1B(256'h8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C),
    .INIT_1C(256'h000000000000000000000000000000000000000000000000A38F8B8C8B8C8C8C),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_5000x8_sub_004096_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(addra[12]),
    .dia({open_n108,open_n109,open_n110,open_n111,open_n112,open_n113,open_n114,open_n115,8'b00000000}),
    .rsta(rsta),
    .doa({open_n137,open_n138,open_n139,open_n140,open_n141,open_n142,open_n143,open_n144,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped),
    .o(doa[7]));

endmodule 

