// Verilog netlist created by TD v4.6.18154
// Wed Nov 11 23:53:31 2020

`timescale 1ns / 1ps
module Bird_Fly  // al_ip/birdfly.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [11:0] addra;  // al_ip/birdfly.v(18)
  input clka;  // al_ip/birdfly.v(19)
  input rsta;  // al_ip/birdfly.v(20)
  output [23:0] doa;  // al_ip/birdfly.v(16)


  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=3600;width=8;num_section=1;width_per_section=8;section_size=24;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSAMUX("1"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFE6E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7878E6FFFFFFFFFFFFE6E6E6E6E6FFFFFF),
    .INIT_0A(256'hE6E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000078E6FFFFFFFFFF7878787878),
    .INIT_0C(256'h0000007878E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFE6E6E6E6E6E6FFFFFFFFE6E6E6FFFFE6E6E6FFE6E6000078E6FFFFFFFF0000),
    .INIT_0E(256'hFF000078E6FF000078FFFFFFFFFFE6E6E6E6FFFFFFFFE6E6FFE6E6E6FFFFFFFF),
    .INIT_0F(256'hE6FFFFFF787878787878E6E6FFFF787878FFE6787878FF7878E6000078E6FFFF),
    .INIT_10(256'h78E6FFFFFF000078E6FFFF00FFFFFFFFFF78787878E6E6FFFF7878E6787878E6),
    .INIT_11(256'h00007878E6E6FF0000000000007878FFFF000000FF78000000FF000078E60000),
    .INIT_12(256'h78E6000078E6FFFFFF000078E6E6FFFFFFFFFFFF000000007878E6E600007800),
    .INIT_13(256'h000000E6FF00007878E6000078E6E6E60000FFFF000078E600000078E6000000),
    .INIT_14(256'hE6FF000078E6000078E6FFFFFF00007878E6E6FFFFFFFF0000E6FF00007878E6),
    .INIT_15(256'h000078E6000078E6FFFF000078E6000078787878E6E6E6FF000078E6FF000078),
    .INIT_16(256'hFF000078E6FF000078E6000078E6FFFFFFFF00007878E6E6FFFF000078E6E6E6),
    .INIT_17(256'h78787878000078E6000078E6FFFF000078E60000000000787878E6E6000078E6),
    .INIT_18(256'h000078E6FF000078E6FF000078E6000078E6FFFFFFFFFF00007878E6E6FF0000),
    .INIT_19(256'hE6E6000000000000000078E6000078E6FFFF000078E6000078E60000007878E6),
    .INIT_1A(256'h000078E6000078E6FF000078E6FF000078E6000078E6FFFFFFFFFFFF00007878),
    .INIT_1B(256'hFF00007878E6FFFFE6E6FFFF000078FF000078E6E6FD000078FD000078E6FFFF),
    .INIT_1C(256'h78FFE6E6000078FF000078E6FF000078E6FF000078E6000078E6FFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFE6E6E6000078E6FF7878E6E6E60000FFFF00007878FFE60000FFFB0000),
    .INIT_1E(256'h55540000547878780000FFFF000078FFFF000078FFFF000078FF000078FFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFF78787878000078FF00007878780000FFFFFF000000E678000055),
    .INIT_20(256'h000057555200005A0000000000FFFEFE0000FFFFFF0000FFFFFF0000FFFF0000),
    .INIT_21(256'hFFFFFFFFFFFFFFFFFF00000000000000FFFFFF0000000000FFFFFFFE00007800),
    .INIT_22(256'h000078E6E6DDDD91E6E66864676271737A7A7677FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE),
    .INIT_24(256'hFFFDFDFE00007878E6E6E678784558555754614F55525554FEFFFFFEFFFEFFFF),
    .INIT_25(256'hFDFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_26(256'hFFFFFFFFFFFFFFFF5500007878780000564556505755604B504F4B52FEFDFCFD),
    .INIT_27(256'h4D5896FDFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_28(256'hFFFFFFFFFFFFFFFFFE675556FFFC0000000000FDFBFF52594A4442585559525E),
    .INIT_29(256'h56525761515695FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFE6A5555FFFEFEFFFFFFFFFFFDFD53544B403E55),
    .INIT_2B(256'h513F443F41495455615F707369FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF7171D4E2E29498E4FEFFFFFDF1E4E05557),
    .INIT_2D(256'hDDDF54554D414246454A54525952585257FDFFFFFFFDFFFFFFFFFFFFFFFFFFFF),
    .INIT_2E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5455EAFDFF5555D4FDFFFFFFEB),
    .INIT_2F(256'hFFFFFCE9DCE055544F474140424F5C5658565D534EFFFFFEFFFFFFFFFFFFFFFF),
    .INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5455EAFDFF5555D4FD),
    .INIT_31(256'h5254D4FDFFFFFFF0DFDF51554E42424743414042423F4144455454C0FFFFFFFF),
    .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5455EAFDFF),
    .INIT_33(256'h55EAFFFF5453D5FDFFFEFEE7D8DD5658504340414443434142454044485455C0),
    .INIT_34(256'h455555C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF54),
    .INIT_35(256'hFFFFFF5455EAFFFFD5D5F4FDFDE5E5B18C804D4D444546444444434343424542),
    .INIT_36(256'h44434844455755C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_37(256'hFFFFFFFFFFFEFF5757E9FCFBFDFFFFFFFFDEE090534C44444242404144444344),
    .INIT_38(256'h4949494949474B4B4D5155C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_39(256'hFFFFFFFFFFFFFFFFF7F7F85554EAFFFFFFFFFFFFFFDDDE834D4B42414444424D),
    .INIT_3A(256'h4442494C5252525252535451505C54C1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFEFF5554545555555454545556565656565143464243),
    .INIT_3C(256'h453E443E454046515454555555555554545455BFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFF56545454555556565555545454545451),
    .INIT_3E(256'h272627394B4645414A494AC3C6D0DDDDDDDDDEDEE1C1C2917877FFFFFFFFFFFF),
    .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF37778322825282725252625252626),
    .INIT_40(256'h000000000000002D57514644505455DCDEEEFFFFFFFFFFFEFFDCDD865553FFFF),
    .INIT_41(256'h5553FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFF154562102000200000000),
    .INIT_42(256'h090909090909090909090822434044464D5055DCE1EFFFFFFFFFFFFFFFDEDD85),
    .INIT_43(256'hFFFFFF935553FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF054541C0A070B),
    .INIT_44(256'h5850525555545454545454545454512A000956564B3C425754BEFFFFFFFFFFFF),
    .INIT_45(256'hFFFFFFFFFFFFFF935553FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_46(256'hFFFFFFFF5659595553545555545554545554542600065650453E445455BEFFFF),
    .INIT_47(256'h4760716FE1E3EEFFFFFFFF955554FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_48(256'hFFFFFFFFFFFFFFFF5551431B1A1B1B1B1B1B1B1B1B1B192A38354746413E4046),
    .INIT_49(256'h3E3E3E3E3C4A5553DFDDEAFFFFFFFF955453FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_4A(256'hFFFFFFFFFFFFFFFFFFFFFFFF5455420003010101010101010101002852523D3E),
    .INIT_4B(256'h554B3C3E3E3E3E3E3E495554E1DFECFFFFFFFF935251FFFFFFFFFFFFFFFFFFFF),
    .INIT_4C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55523E0C0D0B0B0B0B0B0B0B0B0B0B2E),
    .INIT_4D(256'h5555584A3E3B403E3E3E3E3E3E49555455555555555555C0FFFFFFFFFFFFFFFF),
    .INIT_4E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFEFF555255555555555555),
    .INIT_4F(256'h5454545454545648423E3E3E3E3E3E3E3E49555555555555555556BFFEFEFFFF),
    .INIT_50(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF5854545454),
    .INIT_51(256'hD3D4D4D4D4D4D4D4D4D4D36E50505051515151515192D4D4D4D4D4D4D4D4D4EE),
    .INIT_52(256'hFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD4),
    .INIT_53(256'hFFFFFEFEFEFFFFFFFFFFFFFFFFFFFF78555556555555555556A9FFFFFFFFFFFF),
    .INIT_54(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_55(256'hFFFFFFFFFFFFFEFEFFFFFFFFFFFFFFFFFFFFFF78545555555455545455AAFFFF),
    .INIT_56(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_57(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFEFEFFFFFFFFFFFFFF),
    .INIT_58(256'hFFFFFFFFFDFBFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_59(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDFF),
    .INIT_5A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_60(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_61(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_62(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_63(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_64(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_65(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_66(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_67(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_68(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_69(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_70(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_000000_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .dia({open_n52,open_n53,open_n54,open_n55,open_n56,open_n57,open_n58,open_n59,8'b00000000}),
    .rsta(rsta),
    .doa({open_n81,open_n82,open_n83,open_n84,open_n85,open_n86,open_n87,open_n88,doa[7:0]}));
  // address_offset=0;data_offset=8;depth=3600;width=8;num_section=1;width_per_section=8;section_size=24;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSAMUX("1"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFE6E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7878E6FFFFFFFFFFFFE6E6E6E6E6FFFFFF),
    .INIT_0A(256'hE6E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000078E6FFFFFFFFFF7878787878),
    .INIT_0C(256'h0000007878E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFE6E6E6E6E6E6FFFFFFFFE6E6E6FFFFE6E6E6FFE6E6000078E6FFFFFFFF0000),
    .INIT_0E(256'hFF000078E6FF000078FFFFFFFFFFE6E6E6E6FFFFFFFFE6E6FFE6E6E6FFFFFFFF),
    .INIT_0F(256'hE6FFFFFF787878787878E6E6FFFF787878FFE6787878FF7878E6000078E6FFFF),
    .INIT_10(256'h78E6FFFFFF000078E6FFFF00FFFFFFFFFF78787878E6E6FFFF7878E6787878E6),
    .INIT_11(256'h00007878E6E6FF0000000000007878FFFF000000FF78000000FF000078E60000),
    .INIT_12(256'h78E6000078E6FFFFFF000078E6E6FFFFFFFFFFFF000000007878E6E600007800),
    .INIT_13(256'h000000E6FF00007878E6000078E6E6E60000FFFF000078E600000078E6000000),
    .INIT_14(256'hE6FF000078E6000078E6FFFFFF00007878E6E6FFFFFFFF0000E6FF00007878E6),
    .INIT_15(256'h000078E6000078E6FFFF000078E6000078787878E6E6E6FF000078E6FF000078),
    .INIT_16(256'hFF000078E6FF000078E6000078E6FFFFFFFF00007878E6E6FFFF000078E6E6E6),
    .INIT_17(256'h78787878000078E6000078E6FFFF000078E60000000000787878E6E6000078E6),
    .INIT_18(256'h000078E6FF000078E6FF000078E6000078E6FFFFFFFFFF00007878E6E6FF0000),
    .INIT_19(256'hE6E6000000000000000078E6000078E6FFFF000078E6000078E60000007878E6),
    .INIT_1A(256'h000078E6000078E6FF000078E6FF000078E6000078E6FFFFFFFFFFFF00007878),
    .INIT_1B(256'hFF00007878E6FFFFE6E6FFFF000078FF000078E6E6FF000078FF000078E6FEFF),
    .INIT_1C(256'h78FDE6E6000078FF000078E6FF000078E6FF000078E6000078E6FFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFE6E6E6000078E6FF7878E6E6E60000FFFF00007878FDE60000FEFF0000),
    .INIT_1E(256'h494A00004A7878780000FFFF000078FFFF000078FFFF000078FF000078FFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFF78787878000078FF00007878780000FFFFFF000000E67800004A),
    .INIT_20(256'h0000474A4B00004A0000000000FEFEFE0000FFFFFF0000FFFFFF0000FFFF0000),
    .INIT_21(256'hFFFFFFFFFFFFFFFFFF00000000000000FFFFFF0000000000FFFEFFFF00007800),
    .INIT_22(256'h000078E6E6D9DA82E6E6ADAFAEB0AB7271717073FDFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC),
    .INIT_24(256'hFFFFFFFB00007878E6E6E6787852D9D8D9D8D34E494B484BFCFEFEFFFDFFFFFF),
    .INIT_25(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_26(256'hFFFFFEFEFEFEFCFD4C000078787800004855D6D9D8D8D4554D4E4D4FFEFFFCFF),
    .INIT_27(256'h4F498DFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_28(256'hFFFFFFFFFFFFFFFFFF60484BFEFD0000000000FFFEFD4B4892A9A6D7D8D8D8D0),
    .INIT_29(256'hDBDAD7D2504A8DFEFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2A(256'hFFFFFFFFFFFFFFFFFEFFFFFEFD61494AFEFFFDFFFFFFFFFEFFFE494B8EA9AADA),
    .INIT_2B(256'h8DACA9AFB1C3D9D6B8B698686CFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC6A69CFE0DF8D91E1FFFFFEFFEDE4E34A4A),
    .INIT_2D(256'hDDDB49498FABAAA7ABC0D8D8D9DB9F4949FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFD4A4AE7FFFE4949D1FFFEFFFEEC),
    .INIT_2F(256'hFEFFFFEBDDDD4B4A8EA7A9ACA9C1DAD9D9DDA4524FFCFCFCFFFFFFFFFFFFFFFF),
    .INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFD4A4AE9FFFE4949D0FF),
    .INIT_31(256'h4749D0FFFEFFFFECD9DC474A8EA9AAA8A9A9A9A9AAA9A6A7A74A4BBBFFFFFFFF),
    .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFD4A4AE8FFFD),
    .INIT_33(256'h4AE7FEFE4A49D2FFFEFFFCEBDFDB4A4990A9A9AAA9A9A9A9A9A9AAAAAB4849BA),
    .INIT_34(256'hAA4849BBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFD4A),
    .INIT_35(256'hFFFEFD4A4AE8FFFFD0CFF3FFFCE6E7A883878D8CA2AAA9A9A9A9A9A9A9A9AAA9),
    .INIT_36(256'hA9A9A9A8AC4649BBFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_37(256'hFFFFFFFFFFFEFC4B4BE7FEFFFFFFFFFFFFDDDD854855A9A9ABABA8A9AAAAAAAA),
    .INIT_38(256'h9E9F9F9E9F9F9D9EA04849BBFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_39(256'hFFFFFFFFFFFFFFFFF7F6F64B49E5FEFDFDFEFEFEFEDADC8D5963ABABA9A8A9A1),
    .INIT_3A(256'hAAABA1534D4E4E4E4E4D4E4F4F4848BCFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFEFF4C494B4949494B4B4B4A4A4A4A4A4B86A6A8A9AA),
    .INIT_3C(256'hA8AAA7ABA8A8A04C48494A494949494A4A4A4ABAFEFEFFFFFFFFFFFFFFFFFFFF),
    .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE4E4649494948474949494A4A4A4A4A87),
    .INIT_3E(256'h2F2F305A777EACAA8C7774BFBFCAD8D8D8D9D7D6D9BCBB8C7373FFFFFFFFFFFF),
    .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF272733A312F2E2F303030302F2F2F),
    .INIT_40(256'h181818181818182F4852AAA96E4A4BDDDEEEFFFFFEFFFFFEFFDCDD814949FFFF),
    .INIT_41(256'h4949FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE4A4A2C18191517181818),
    .INIT_42(256'h1C1C1C1C1C1C1C1C1C1C1D2E3E4DA2A3725152DEDCEDFFFFFEFFFFFFFFDEDD80),
    .INIT_43(256'hFFFFFF8E4949FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE4A4A2C1C1C1D),
    .INIT_44(256'h4B4C4B494A4A4A4A4A4A4A4A4A4A4A2E191D4B4A738A844E4AB9FEFFFFFFFFFF),
    .INIT_45(256'hFEFFFFFFFFFFFF8E4949FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFEFE),
    .INIT_46(256'hFFFFFFFF4B494747494747474747474747474630191C494A7487804F4BBBFFFF),
    .INIT_47(256'h76726969E1E1EDFFFFFFFF8E4949FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_48(256'hFFFFFFFFFFFFFFFF4B4B40282A282828282828282828272E383F757882888679),
    .INIT_49(256'h878787878868494ADCDDEAFFFFFFFF8E494AFEFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_4A(256'hFFFFFFFFFFFFFFFFFFFFFFFF4B4939181817171717171717171719304B518687),
    .INIT_4B(256'h50588687878787878768494ADADCE9FEFEFEFD8F4B4CFEFFFFFFFFFFFFFFFFFF),
    .INIT_4C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4B4A3E1E201F1F1F1F1F1F1F1F1F2036),
    .INIT_4D(256'h4949466A888888878787878788684A4A4A49494949494BBAFEFFFFFFFFFFFFFF),
    .INIT_4E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFE4A4949494949494949),
    .INIT_4F(256'h4A4A4A4A4A4A486A878787878787878788674A494949494949494ABAFEFFFFFF),
    .INIT_50(256'hFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFD4B494A4A4A),
    .INIT_51(256'hD1D1D1D1D1D1D1D1D1D1D16F56565655555555555593D1D1D1D1D1D1D1D1D1ED),
    .INIT_52(256'hFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFED1),
    .INIT_53(256'hFFFFFDFEFEFFFFFFFFFFFFFFFFFFFE704949494A4A4A4A4A4AA3FEFFFFFFFFFF),
    .INIT_54(256'hFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_55(256'hFFFFFFFFFFFFFEFEFFFFFFFFFFFFFFFFFFFFFE7149494A494A494A4A49A4FFFF),
    .INIT_56(256'hFDFEFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_57(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFDFFFFFFFFFFFFFF),
    .INIT_58(256'hFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_59(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFEFFFFFE),
    .INIT_5A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_60(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_61(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_62(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_63(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_64(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_65(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_66(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_67(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_68(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_69(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_70(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_000000_008 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .dia({open_n110,open_n111,open_n112,open_n113,open_n114,open_n115,open_n116,open_n117,8'b00000000}),
    .rsta(rsta),
    .doa({open_n139,open_n140,open_n141,open_n142,open_n143,open_n144,open_n145,open_n146,doa[15:8]}));
  // address_offset=0;data_offset=16;depth=3600;width=8;num_section=1;width_per_section=8;section_size=24;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSAMUX("1"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7878FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000078FFFFFFFFFFFF7878787878),
    .INIT_0C(256'h0000007878FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000078FFFFFFFFFF0000),
    .INIT_0E(256'hFF000078FFFF000078FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFF787878787878FFFFFFFF787878FFFF787878FF7878FF000078FFFFFF),
    .INIT_10(256'h78FFFFFFFF000078FFFFFF00FFFFFFFFFF78787878FFFFFFFF7878FF787878FF),
    .INIT_11(256'h00007878FFFFFF0000000000007878FFFF000000FF78000000FF000078FF0000),
    .INIT_12(256'h78FF000078FFFFFFFF000078FFFFFFFFFFFFFFFF000000007878FFFF00007800),
    .INIT_13(256'h000000FFFF00007878FF000078FFFFFF0000FFFF000078FF00000078FF000000),
    .INIT_14(256'hFFFF000078FF000078FFFFFFFF00007878FFFFFFFFFFFF0000FFFF00007878FF),
    .INIT_15(256'h000078FF000078FFFFFF000078FF000078787878FFFFFFFF000078FFFF000078),
    .INIT_16(256'hFF000078FFFF000078FF000078FFFFFFFFFF00007878FFFFFFFF000078FFFFFF),
    .INIT_17(256'h78787878000078FF000078FFFFFF000078FF0000000000787878FFFF000078FF),
    .INIT_18(256'h000078FFFF000078FFFF000078FF000078FFFFFFFFFFFF00007878FFFFFF0000),
    .INIT_19(256'hFFFF000000000000000078FF000078FFFFFF000078FF000078FF0000007878FF),
    .INIT_1A(256'h000078FF000078FFFF000078FFFF000078FF000078FFFFFFFFFFFFFF00007878),
    .INIT_1B(256'hFF00007878FFFFFFFFFFFFFF000078FF000078FFFFFE000078FF000078FFFFFC),
    .INIT_1C(256'h78FFFFFF000078FF000078FFFF000078FFFF000078FF000078FFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFF000078FFFF7878FFFFFF0000FFFF00007878FFFF0000FFFF0000),
    .INIT_1E(256'h5C5B00005B7878780000FFFF000078FFFF000078FFFF000078FF000078FFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFF78787878000078FF00007878780000FFFFFF000000FF7800005A),
    .INIT_20(256'h00005E5B5500005C0000000000FFFFFE0000FFFFFF0000FFFFFF0000FFFF0000),
    .INIT_21(256'hFFFFFFFFFFFFFFFFFF00000000000000FFFFFF0000000000FFFFFFFD00007800),
    .INIT_22(256'h000078FFFFDEDE95FFFF65696A676F757D7D7B79FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_24(256'hFEFEFFFF00007878FFFFFF78784D5459585A5E565D595B59FFFFFDFBFFFCFFFF),
    .INIT_25(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_26(256'hFEFFFFFFFFFFFFFF590000787878000060485A57575B5D4C55545450FEFEFFFF),
    .INIT_27(256'h545A9BFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_28(256'hFFFFFFFFFFFFFFFFFE695E59FFFE0000000000FFFDFF5B5E2102085557565665),
    .INIT_29(256'h59555A63545B98FFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2A(256'hFFFFFFFFFFFFFFFFFFFFFFFEFD6C5E58FEFEFEFFFFFFFCFFFDFF5D5826050256),
    .INIT_2B(256'h270102161837535865656F7671FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF7474D5E3E3969AE4FDFFFFFFF2DDE7585A),
    .INIT_2D(256'hDDE05C5B25010106032C585A54595D5E5AFEFEFFFEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_2E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5B5AEBFFFF5B5DD6FFFFFFFFE9),
    .INIT_2F(256'hFFFEFCEBDDDC595B24060300042B52565552524B50FFFFFEFFFFFFFFFFFFFFFF),
    .INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5B5AEBFFFF5B5BD6FF),
    .INIT_31(256'h585BD6FFFFFEFEEDE3DD5C59240002030304050403050806085958C3FFFFFFFF),
    .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5B5AEBFFFF),
    .INIT_33(256'h5AEBFFFF5A59D6FFFFFDFFE8D9E1595E240406030303030403030300005E5BC4),
    .INIT_34(256'h005E5BC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5B),
    .INIT_35(256'hFFFFFF5B5AEBFFFDD6D6F4FEFEE5E3B2898020200D0103030202030303030204),
    .INIT_36(256'h0203010501605DC2FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_37(256'hFFFFFFFFFEFFFF5D5AEAFCFFFFFDFFFEFFDDDC905C4804020001030401010101),
    .INIT_38(256'h171616171616171817585DC2FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_39(256'hFFFFFFFFFFFFFFFFF8F9F85C5AEAFFFFFFFFFFFFFFDEE2804634020104060214),
    .INIT_3A(256'h01030E4A5353535353545350555C5CC3FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFEFF585B585B5B5B5959595A5A5A5A5A5A2D0C060302),
    .INIT_3C(256'h0303040304040D515A5A5B5B5B5B5B585B5A5BC1FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF555D5D5D5B5E5E5D5D5D5B5B5B5B602D),
    .INIT_3E(256'hBDBDBE722A2401041A2C33BFC9D3E0E1E0E0E1E1DFC4C5967A7CFFFFFFFFFFFF),
    .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF47A7AA0BCBDBDBBBBBBBBBBBDBDBD),
    .INIT_40(256'hFEFEFEFEFEFEFEAC5B4C0204385959DEDDEDFEFFFFFFFFFEFFDCDD8B5B5BFFFF),
    .INIT_41(256'h5B5BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF15C5CCCF9FDFFFFFEFEFE),
    .INIT_42(256'hF1F2F2F2F2F2F2F2F2F2F3B2775F0F0E314E4FDFE0EEFFFFFFFFFFFFFFDEDD8A),
    .INIT_43(256'hFFFFFF975B5BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF1595ABFF3F2F0),
    .INIT_44(256'h58575A5D595A5B5A5A5B5A5A5B5A59BDFCF05859290B12555AC0FFFFFFFFFFFF),
    .INIT_45(256'hFFFFFFFFFFFFFF975B5BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_46(256'hFFFFFEFF575B5D5E5D5F5F5F5F5F5F5F5F5F60BCFFF35C58290E175257BFFFFF),
    .INIT_47(256'h274F7473E1E1EDFFFFFFFF975D59FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_48(256'hFFFFFFFFFFFFFFFF585877CFCFD0D0D0D0D0D0D0D0D0D4B28E802523150A0E23),
    .INIT_49(256'h0B0B0B0B0B335B5ADEDDEAFFFFFFFF975D59FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_4A(256'hFFFFFFFFFFFFFFFFFFFFFFFF595C83FEFEFFFFFFFFFFFFFFFFFFFBAD5A4B0A0B),
    .INIT_4B(256'h4D410C0B0B0B0B0B0B335B5AE1DDEBFEFEFFFF975956FFFFFFFFFFFFFFFFFFFF),
    .INIT_4C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF575A7BEDEBEBEBEBEBEBEBEBEBEBEB9D),
    .INIT_4D(256'h5B5B5D330B0B090B0B0B0B0B0A335A5B5A5B5B5B5B5D5BC4FFFEFFFFFFFFFFFF),
    .INIT_4E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFEFF5D5B5B5B5B5B5B5B5B),
    .INIT_4F(256'h5A5A5A5A5A5A5A330A0B0B0B0B0B0B0B0A355A5D5D5B5B5B5B5B5DC3FEFEFFFF),
    .INIT_50(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFF5D595A5A5A),
    .INIT_51(256'hD4D5D5D5D5D5D5D5D5D5D46C4A48494A4A4A4A4A4B90D4D5D5D5D5D5D5D5D5EF),
    .INIT_52(256'hFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD5),
    .INIT_53(256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFF7B5B5C5C5A5A5A5A5A5DAAFFFFFFFFFFFF),
    .INIT_54(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_55(256'hFFFFFFFFFFFFFEFEFFFFFFFFFFFFFFFFFFFFFE785A5A595B5B5B5B5B5AABFEFE),
    .INIT_56(256'hFEFEFEFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_57(256'hFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFDFEFFFFFEFFFFFFFFFF),
    .INIT_58(256'hFFFFFFFFFEFDFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_59(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFDFEFEFFFF),
    .INIT_5A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_5F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_60(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_61(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_62(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_63(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_64(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_65(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_66(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_67(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_68(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_69(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_6F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_70(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_000000_016 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .dia({open_n168,open_n169,open_n170,open_n171,open_n172,open_n173,open_n174,open_n175,8'b00000000}),
    .rsta(rsta),
    .doa({open_n197,open_n198,open_n199,open_n200,open_n201,open_n202,open_n203,open_n204,doa[23:16]}));

endmodule 

