// Verilog netlist created by TD v4.6.18154
// Sat Nov  7 11:31:16 2020

`timescale 1ns / 1ps
module Bird_Fly  // ../Bin/AngryBird_Demo/al_ip/birdggg.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [11:0] addra;  // ../Bin/AngryBird_Demo/al_ip/birdggg.v(18)
  input clka;  // ../Bin/AngryBird_Demo/al_ip/birdggg.v(19)
  input rsta;  // ../Bin/AngryBird_Demo/al_ip/birdggg.v(20)
  output [23:0] doa;  // ../Bin/AngryBird_Demo/al_ip/birdggg.v(16)

  wire [0:1] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b10/B0_0 ;
  wire  \inst_doa_mux_b10/B0_1 ;
  wire  \inst_doa_mux_b11/B0_0 ;
  wire  \inst_doa_mux_b11/B0_1 ;
  wire  \inst_doa_mux_b12/B0_0 ;
  wire  \inst_doa_mux_b12/B0_1 ;
  wire  \inst_doa_mux_b13/B0_0 ;
  wire  \inst_doa_mux_b13/B0_1 ;
  wire  \inst_doa_mux_b14/B0_0 ;
  wire  \inst_doa_mux_b14/B0_1 ;
  wire  \inst_doa_mux_b15/B0_0 ;
  wire  \inst_doa_mux_b15/B0_1 ;
  wire  \inst_doa_mux_b16/B0_0 ;
  wire  \inst_doa_mux_b16/B0_1 ;
  wire  \inst_doa_mux_b17/B0_0 ;
  wire  \inst_doa_mux_b17/B0_1 ;
  wire  \inst_doa_mux_b18/B0_0 ;
  wire  \inst_doa_mux_b18/B0_1 ;
  wire  \inst_doa_mux_b19/B0_0 ;
  wire  \inst_doa_mux_b19/B0_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b20/B0_0 ;
  wire  \inst_doa_mux_b20/B0_1 ;
  wire  \inst_doa_mux_b21/B0_0 ;
  wire  \inst_doa_mux_b21/B0_1 ;
  wire  \inst_doa_mux_b22/B0_0 ;
  wire  \inst_doa_mux_b22/B0_1 ;
  wire  \inst_doa_mux_b23/B0_0 ;
  wire  \inst_doa_mux_b23/B0_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b9/B0_0 ;
  wire  \inst_doa_mux_b9/B0_1 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i0_011;
  wire inst_doa_i0_012;
  wire inst_doa_i0_013;
  wire inst_doa_i0_014;
  wire inst_doa_i0_015;
  wire inst_doa_i0_016;
  wire inst_doa_i0_017;
  wire inst_doa_i0_018;
  wire inst_doa_i0_019;
  wire inst_doa_i0_020;
  wire inst_doa_i0_021;
  wire inst_doa_i0_022;
  wire inst_doa_i0_023;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i1_009;
  wire inst_doa_i1_010;
  wire inst_doa_i1_011;
  wire inst_doa_i1_012;
  wire inst_doa_i1_013;
  wire inst_doa_i1_014;
  wire inst_doa_i1_015;
  wire inst_doa_i1_016;
  wire inst_doa_i1_017;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i2_009;
  wire inst_doa_i2_010;
  wire inst_doa_i2_011;
  wire inst_doa_i2_012;
  wire inst_doa_i2_013;
  wire inst_doa_i2_014;
  wire inst_doa_i2_015;
  wire inst_doa_i2_016;
  wire inst_doa_i2_017;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;
  wire inst_doa_i3_008;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[10]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[11]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'h700C4203847C3C8F81E3103C03FFFFFFFFFFC3E03FFFFFFFFFFE3F07FFFFFFFF),
    .INITP_02(256'h000C00008403C0C000C0010840381E20080030000383F00002018840386F8180),
    .INITP_03(256'hFC04070080318C47E02030844108403F83310441008403F00000C00008403E04),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFE6E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7878E6FFFFFFFFFFFFE6E6E6E6E6FFFFFF),
    .INIT_0A(256'hE6E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000078E6FFFFFFFFFF7878787878),
    .INIT_0C(256'h0000007878E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFE6E6E6E6E6E6FFFFFFFFE6E6E6FFFFE6E6E6FFE6E6000078E6FFFFFFFF0000),
    .INIT_0E(256'hFF000078E6FF000078FFFFFFFFFFE6E6E6E6FFFFFFFFE6E6FFE6E6E6FFFFFFFF),
    .INIT_0F(256'hE6FFFFFF787878787878E6E6FFFF787878FFE6787878FF7878E6000078E6FFFF),
    .INIT_10(256'h78E6FFFFFF000078E6FFFF00FFFFFFFFFF78787878E6E6FFFF7878E6787878E6),
    .INIT_11(256'h00007878E6E6FF0000000000007878FFFF000000FF78000000FF000078E60000),
    .INIT_12(256'h78E6000078E6FFFFFF000078E6E6FFFFFFFFFFFF000000007878E6E600007800),
    .INIT_13(256'h000000E6FF00007878E6000078E6E6E60000FFFF000078E600000078E6000000),
    .INIT_14(256'hE6FF000078E6000078E6FFFFFF00007878E6E6FFFFFFFF0000E6FF00007878E6),
    .INIT_15(256'h000078E6000078E6FFFF000078E6000078787878E6E6E6FF000078E6FF000078),
    .INIT_16(256'hFF000078E6FF000078E6000078E6FFFFFFFF00007878E6E6FFFF000078E6E6E6),
    .INIT_17(256'h78787878000078E6000078E6FFFF000078E60000000000787878E6E6000078E6),
    .INIT_18(256'h000078E6FF000078E6FF000078E6000078E6FFFFFFFFFF00007878E6E6FF0000),
    .INIT_19(256'hE6E6000000000000000078E6000078E6FFFF000078E6000078E60000007878E6),
    .INIT_1A(256'h000078E6000078E6FF000078E6FF000078E6000078E6FFFFFFFFFFFF00007878),
    .INIT_1B(256'hFF00007878E6FFFFE6E6FFFF000078FF000078E6E6FD000078FD000078E6FFFF),
    .INIT_1C(256'h78FFE6E6000078FF000078E6FF000078E6FF000078E6000078E6FFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFE6E6E6000078E6FF7878E6E6E60000FFFF00007878FFE60000FFFB0000),
    .INIT_1E(256'h55540000547878780000FFFF000078FFFF000078FFFF000078FF000078FFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFF78787878000078FF00007878780000FFFFFF000000E678000055),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n63,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_008,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hF03C62478C7FFFFFFFFFFC7C07FFFFFFFFFFC7E0FFFFFFFFFFFE7FFFFFFFFFFF),
    .INITP_02(256'h011C40318C47C3C711C40F18C4787E6118473108478FF0300E01884478EF8791),
    .INITP_03(256'hFC04071148318C47FC6730CC7118C47F87F11C46118C47F0C011C44118C47E1C),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFF3F3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3C3CF3FFFFFFFFFFFFF3F3F3F3F3FFFFFF),
    .INIT_0A(256'hF3F3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00003CF3FFFFFFFFFF3C3C3C3C3C),
    .INIT_0C(256'h0000003C3CF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFF3F3F3F3F3F3FFFFFFFFF3F3F3FFFFF3F3F3FFF3F300003CF3FFFFFFFF0000),
    .INIT_0E(256'hFF00003CF3FF00003CFFFFFFFFFFF3F3F3F3FFFFFFFFF3F3FFF3F3F3FFFFFFFF),
    .INIT_0F(256'hF3FFFFFF3C3C3C3C3C3CF3F3FFFF3C3C3CFFF33C3C3CFF3C3CF300003CF3FFFF),
    .INIT_10(256'h3CF3FFFFFF00003CF3FFFF00FFFFFFFFFF3C3C3C3CF3F3FFFF3C3CF33C3C3CF3),
    .INIT_11(256'h00003C3CF3F3FF0000000000003C3CFFFF000000FF3C000000FF00003CF30000),
    .INIT_12(256'h3CF300003CF3FFFFFF00003CF3F3FFFFFFFFFFFF000000003C3CF3F300003C00),
    .INIT_13(256'h000000F3FF00003C3CF300003CF3F3F30000FFFF00003CF30000003CF3000000),
    .INIT_14(256'hF3FF00003CF300003CF3FFFFFF00003C3CF3F3FFFFFFFF0000F3FF00003C3CF3),
    .INIT_15(256'h00003CF300003CF3FFFF00003CF300003C3C3C3CF3F3F3FF00003CF3FF00003C),
    .INIT_16(256'hFF00003CF3FF00003CF300003CF3FFFFFFFF00003C3CF3F3FFFF00003CF3F3F3),
    .INIT_17(256'h3C3C3C3C00003CF300003CF3FFFF00003CF300000000003C3C3CF3F300003CF3),
    .INIT_18(256'h00003CF3FF00003CF3FF00003CF300003CF3FFFFFFFFFF00003C3CF3F3FF0000),
    .INIT_19(256'hF3F300000000000000003CF300003CF3FFFF00003CF300003CF30000003C3CF3),
    .INIT_1A(256'h00003CF300003CF3FF00003CF3FF00003CF300003CF3FFFFFFFFFFFF00003C3C),
    .INIT_1B(256'hFF00003C3CF3FFFFF3F3FFFF00003CFF00003CF3F37F00003CFF00003CF3FF7F),
    .INIT_1C(256'h3CFEF3F300003CFF00003CF3FF00003CF3FF00003CF300003CF3FFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFF3F3F300003CF3FF3C3CF3F3F30000FFFF00003C3CFEF30000FFFF0000),
    .INIT_1E(256'h24A50000A53C3C3C0000FFFF00003CFFFF00003CFFFF00003CFF00003CFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFF3C3C3C3C00003CFF00003C3C3C0000FFFFFF000000F33C000025),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_000000_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n106,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_017,inst_doa_i0_016,inst_doa_i0_015,inst_doa_i0_014,inst_doa_i0_013,inst_doa_i0_012,inst_doa_i0_011,inst_doa_i0_010,inst_doa_i0_009}));
  // address_offset=0;data_offset=18;depth=3600;width=2;num_section=1;width_per_section=2;section_size=24;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFF0BFFEAAFFFFFFFFFFFFFFFFFFFFFFFEBFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFAAAFFABEAEB0BFC2F0BFFFFFFFFFFFFFFFFFFFFFF0BFF002BFFFFFFFFFFFFF),
    .INIT_04(256'h03C2B0BF0F0B02C0B0BFC2FFFF00AF080AFC002BC0E030B0BFC2FCFFEABFEBAB),
    .INIT_05(256'hAA0B0BF0B002AF0BC2F0B0BFF0AFF0BF0B0BF0B0AAFF0BC2F0B0BFC2BFFC3C2B),
    .INIT_06(256'hC2BFFF0B0BF0B0BF0B0BC2F0B0BFFF0AF0000B0BF0B0B02B0BC2F0B0BFFC2BF0),
    .INIT_07(256'hFFFAA0B0A83F0382E0AA0F0BC2F0B0BFFFF0BEBF0F0AF0F0BF0B0BC2F0B0BFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFF0BFDF69DFAFFFFFFFFFFC000FC00FF080E43003F0FC3F0F0),
    .INIT_09(256'h6BBFFFFFFFFFFFFFFFFF82A0296F54FFFFFFFFFFFFFFFFFFFF0AFEB6ADEAFEFF),
    .INIT_0A(256'h41925D3FFFFFFFFFFFFFFFFEFFFFFE51986BFFFFFFFFFFFFFFFFEEF003FB0955),
    .INIT_0B(256'hFEFA5061423FFFFFFFFFFFFFFEAFB7FECE413A6FBFFFFFFFFFFFFFFD5067FCDA),
    .INIT_0C(256'hAFA7FE8B54010039FFFFFFFFFFFFFEAFA7FF3E401519A8FFFFFFFFFFFFFEAFA7),
    .INIT_0D(256'hFFFFAFFFFCE40100010CFFFFFFFFFFFFFEAF57D080C0000138FFFFFFFFFFFFFE),
    .INIT_0E(256'hFFFFFFAAAAAAABD00E00107CFFFFFFFFFFFFABAFFFF0505155566CFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFDA3FAABFFC91B38000D5BFFFFFFFFFFF7FBFFAA3045CAAAAA8FFFFFF),
    .INIT_10(256'hFDAFFFFFFFFFCAC00000007F3F3FFFFEAFFFFFFFFFCFEFFFFFFFB1ABFFFFFEAF),
    .INIT_11(256'h740FFDEFFFFFFFFFFF6FFFFFF3CEB47FFFFDAFFFFFFFFFFF9BAAAAABCAA18FFF),
    .INIT_12(256'hCEAA8A3BFD9FFFFFFFFFFFB3FFFFFBAAAA8AFBFDEFFFFFFFFFFFA7C00004C46C),
    .INIT_13(256'hAAA8AAAA9BEAACFFFFFFFFFFFFFFAAAAACAAAA8AAAB9FFFFFFFFFFFF6BAAAAAB),
    .INIT_14(256'hFFFFFFFEBEAAEFFFFFFFFFFFFFFFFFFD555557AAAA855557FFFFFFFFFFFFFFAA),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h00000000000000000000000000000000000000000000000000000000FFFFFFFF),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_000000_018 (
    .addra({addra,1'b1}),
    .clka(clka),
    .dia({open_n155,open_n156,open_n157,1'b0,open_n158,open_n159,1'b0,open_n160,open_n161}),
    .rsta(rsta),
    .doa({open_n176,open_n177,open_n178,open_n179,open_n180,open_n181,open_n182,inst_doa_i0_019,inst_doa_i0_018}));
  // address_offset=0;data_offset=20;depth=3600;width=2;num_section=1;width_per_section=2;section_size=24;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFF0FFC3F0FFFFFFFFFFFFFFFFFFFFFFF0FFF003FFFFFFFFFFFFFF),
    .INIT_04(256'h03C3F0FF0F0F03C0F0FFC3FFFF00FF0C0FFC003FC0F030F0FFC3FCFFFFFFFFFF),
    .INIT_05(256'hFF0F0FF0F003FF0FC3F0F0FFF0FFF0FF0F0FF0F0FFFF0FC3F0F0FFC3FFFC3C3F),
    .INIT_06(256'hC3FFFF0F0FF0F0FF0F0FC3F0F0FFFF0FF0000F0FF0F0F03F0FC3F0F0FFFC3FF0),
    .INIT_07(256'hFFFFF0F0FC3F03C1507F0F0FC3F0F0FFFFF0FFFF0F0FF0F0FF0F0FC3F0F0FFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFF0FD5FAABFFFFFFFFFFFFC000FC00FF0C0541003F0FC3F0F0),
    .INIT_09(256'h57FFFFFFFFFFFFFFFFFF43F0855455FFFFFFFFFFFFFFFFFFFF0FFFC55555FFFF),
    .INIT_0A(256'h8175ABFFFFFFFFFFFFFFFFE5FFFFF5815657FFFFFFFFFFFFFFFFE5F003F58156),
    .INIT_0B(256'hFE558025547FFFFFFFFFFFFFFD6F57FE658025557FFFFFFFFFFFFFFFDA5BFF65),
    .INIT_0C(256'h6F57FE6580000014FFFFFFFFFFFFFD6F57FE9580000014FFFFFFFFFFFFFD6F57),
    .INIT_0D(256'hFFFD6FFFD54000000024FFFFFFFFFFFFFD6F5FEB0A00000014FFFFFFFFFFFFFD),
    .INIT_0E(256'hFFFFFF555555560000555554FFFFFFFFFFFFFD6FFFD83001555554FFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFBFFFFFFFA06F1AAA41FFFFFFFFFFFF5555555A0001555554FFFFFF),
    .INIT_10(256'hFD5FFFFFFFFFF5FFFFFFFFD0C1AFFFD45FFFFFFFFFF53FFFFFFE40D56FFFD45F),
    .INIT_11(256'h8FABFD5FFFFFFFFFFF5555555BF5857FFFFD5FFFFFFFFFFF55555557F5854FFF),
    .INIT_12(256'h0000359BFD5FFFFFFFFFFF53FFFFFE4000355BFD5FFFFFFFFFFF5C1555570A42),
    .INIT_13(256'h55570000355554FFFFFFFFFFFFFD5555570000355554FFFFFFFFFFFF5EAAAAA9),
    .INIT_14(256'hFFFFFFFF55556FFFFFFFFFFFFFFFFFFD5555560000155556FFFFFFFFFFFFFD55),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55556FFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h00000000000000000000000000000000000000000000000000000000FFFFFFFF),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_000000_020 (
    .addra({addra,1'b1}),
    .clka(clka),
    .dia({open_n214,open_n215,open_n216,1'b0,open_n217,open_n218,1'b0,open_n219,open_n220}),
    .rsta(rsta),
    .doa({open_n235,open_n236,open_n237,open_n238,open_n239,open_n240,open_n241,inst_doa_i0_021,inst_doa_i0_020}));
  // address_offset=0;data_offset=22;depth=3600;width=2;num_section=1;width_per_section=2;section_size=24;working_depth=4096;working_width=2;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("2"),
    .DATA_WIDTH_B("2"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFF07FFD55FFFFFFFFFFFFFFFFFFFFFFFD7FFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFF555FF57D5D707FC1F07FFFFFFFFFFFFFFFFFFFFFF07FF0017FFFFFFFFFFFFF),
    .INIT_04(256'h03C1707F0F0701C0707FC1FFFF005F0405FC0017C0D030707FC1FCFFD57FD757),
    .INIT_05(256'h550707F070015F07C1F0707FF05FF07F0707F07055FF07C1F0707FC17FFC3C17),
    .INIT_06(256'hC17FFF0707F0707F0707C1F0707FFF05F0000707F070701707C1F0707FFC17F0),
    .INIT_07(256'hFFF55070543F034150550F07C1F0707FFFF07D7F0F05F0F07F0707C1F0707FFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFF07FEF55555FFFFFFFFFFC000FC00FF040541003F0FC3F0F0),
    .INIT_09(256'h5BFFFFFFFFFFFFFFFFFF4150555555FFFFFFFFFFFFFFFFFFFF05FD555555FFFF),
    .INIT_0A(256'h0005557FFFFFFFFFFFFFFFD5FFFFF501555BFFFFFFFFFFFFFFFFD5F003F50155),
    .INIT_0B(256'hFFF50005557FFFFFFFFFFFFFFD7F5FFFF50005557FFFFFFFFFFFFFFD7FAFFFF5),
    .INIT_0C(256'h7F5FFFF500000017FFFFFFFFFFFFFD7F5FFFF500000017FFFFFFFFFFFFFD7F5F),
    .INIT_0D(256'hFFFD7FFFFE5000000017FFFFFFFFFFFFFD7FFFFEA000000017FFFFFFFFFFFFFD),
    .INIT_0E(256'hFFFFFF555555540001555557FFFFFFFFFFFFFD7FFFFE4000000017FFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFF5AAAAAAA90002FFFFFE5FFFFFFFFFFF555555540001555557FFFFFF),
    .INIT_10(256'hFE5FFFFFFFFFF5BFFFFFFE5017FFFFFE5FFFFFFFFFF5FFFFFFFE5017FFFFFE5F),
    .INIT_11(256'h15FFFE5FFFFFFFFFFF55555556F5016FFFFE5FFFFFFFFFFF55555556F5017FFF),
    .INIT_12(256'h500005FFFE5FFFFFFFFFFF5BFFFFFE500005FFFE5FFFFFFFFFFF57FFFFFEA000),
    .INIT_13(256'h55540000055557FFFFFFFFFFFFFD5555540000055557FFFFFFFFFFFF57FFFFFE),
    .INIT_14(256'hFFFFFFFD55556FFFFFFFFFFFFFFFFFFFFFFFFD55556FFFFFFFFFFFFFFFFFFD55),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55556FFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h00000000000000000000000000000000000000000000000000000000FFFFFFFF),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_000000_022 (
    .addra({addra,1'b1}),
    .clka(clka),
    .dia({open_n273,open_n274,open_n275,1'b0,open_n276,open_n277,1'b0,open_n278,open_n279}),
    .rsta(rsta),
    .doa({open_n294,open_n295,open_n296,open_n297,open_n298,open_n299,open_n300,inst_doa_i0_023,inst_doa_i0_022}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFC10051B5FFFFFFFFF002AD1FFFFFFFFE0432DFFFFF80E0B0280039CC),
    .INITP_01(256'h7E6DC8FFFFFFA6F4FD8FFFFFFFFCDFB4BE03FFFFFF6E7EB4A2FFFFFFFF941650),
    .INITP_02(256'hF9DFF7D0E3BFFFFFA372E3FD3FFFFFFA455D6FCAFFFFFFA3D6A4F5BFFFFFFA6D),
    .INITP_03(256'hFFFF9687C8586AFFFFFE3BC1305E03FFFFD7F8227858BFFFFF9D81FB6E3BFFFF),
    .INIT_00(256'h000057555200005A0000000000FFFEFE0000FFFFFF0000FFFFFF0000FFFF0000),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFF00000000000000FFFFFF0000000000FFFFFFFE00007800),
    .INIT_02(256'h000078E6E6DDDD91E6E66864676271737A7A7677FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE),
    .INIT_04(256'hFFFDFDFE00007878E6E6E678784558555754614F55525554FEFFFFFEFFFEFFFF),
    .INIT_05(256'hFDFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFF5500007878780000564556505755604B504F4B52FEFDFCFD),
    .INIT_07(256'h4D5896FDFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFE675556FFFC0000000000FDFBFF52594A4442585559525E),
    .INIT_09(256'h56525761515695FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFE6A5555FFFEFEFFFFFFFFFFFDFD53544B403E55),
    .INIT_0B(256'h513F443F41495455615F707369FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF7171D4E2E29498E4FEFFFFFDF1E4E05557),
    .INIT_0D(256'hDDDF54554D414246454A54525952585257FDFFFFFFFDFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5455EAFDFF5555D4FDFFFFFFEB),
    .INIT_0F(256'hFFFFFCE9DCE055544F474140424F5C5658565D534EFFFFFEFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5455EAFDFF5555D4FD),
    .INIT_11(256'h5254D4FDFFFFFFF0DFDF51554E42424743414042423F4144455454C0FFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5455EAFDFF),
    .INIT_13(256'h55EAFFFF5453D5FDFFFEFEE7D8DD5658504340414443434142454044485455C0),
    .INIT_14(256'h455555C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF54),
    .INIT_15(256'hFFFFFF5455EAFFFFD5D5F4FDFDE5E5B18C804D4D444546444444434343424542),
    .INIT_16(256'h44434844455755C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFEFF5757E9FCFBFDFFFFFFFFDEE090534C44444242404144444344),
    .INIT_18(256'h4949494949474B4B4D5155C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFF7F7F85554EAFFFFFFFFFFFFFFDDDE834D4B42414444424D),
    .INIT_1A(256'h4442494C5252525252535451505C54C1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFEFF5554545555555454545556565656565143464243),
    .INIT_1C(256'h453E443E454046515454555555555554545455BFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFF56545454555556565555545454545451),
    .INIT_1E(256'h272627394B4645414A494AC3C6D0DDDDDDDDDEDEE1C1C2917877FFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF37778322825282725252625252626),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n326,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_008,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  // address_offset=1024;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h7FFFFFFFFF003C0FFFFFFFFFF0E072DBFFFFFFFF1ECE2FFFFF80E0E0300739CC),
    .INITP_01(256'hD16777FFFFFFFFBE1191FFFFFFFE3CF5B637FFFFFFF2FD4B35FFFFFFFFAC174E),
    .INITP_02(256'hFEDB8120C1FFFFFFFEDB03FE7FFFFFFFFBA13EE6FFFFFFFF7E83891FFFFFFFFF),
    .INITP_03(256'hFFFFB0F838B409BFFFFF0E3CD0FEEFFFFFF5C7E77FA1FFFFFF0FFEA6FE9FFFFF),
    .INIT_00(256'h000023A5A50000250000000000FFFF7F0000FFFFFF0000FFFFFF0000FFFF0000),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFF00000000000000FFFFFF0000000000FFFFFFFF00003C00),
    .INIT_02(256'h00003CF3F36C6DC1F3F3D6D757D8D5B9B8B8B8B9FEFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE),
    .INIT_04(256'h7F7FFFFD00003C3CF3F3F33C3CA96CEC6C6C6927A4A5A4A5FEFFFFFFFE7FFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'h7FFFFFFFFFFFFEFEA600003C3C3C0000242A6BECECECEA2AA62726277F7FFEFF),
    .INIT_07(256'h2724C6FF7FFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFF7FB024A5FF7E0000000000FFFFFEA524C95453EBEC6C6CE8),
    .INIT_09(256'hEDED6BE928A546FFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFF7FFE3024257F7F7EFFFFFF7FFFFFFFA42547D4556D),
    .INIT_0B(256'hC6D6545758E1EC6BDCDBCC34B67EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFF7FFFFE3534E7F0EF464870FFFFFFFF76F2F12525),
    .INIT_0D(256'hEE6D24A4C7D5D553D5606C6C6CEDCF24247F7FFF7FFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA525F3FFFFA4A468FFFFFFFFF6),
    .INIT_0F(256'hFF7F7FF5EE6EA5A54753D45654E06D6CEC6E52A927FEFE7EFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA525F4FFFFA4A468FF),
    .INIT_11(256'h23A468FFFF7F7FF6ECEE23A5475455D4D454D454D5D4535353A525DDFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA525F4FFFE),
    .INIT_13(256'h25F3FFFF25A469FFFFFFFE75EFEDA524485454D5D4D4D454D4D4D5555524A45D),
    .INIT_14(256'h5524A4DDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA5),
    .INIT_15(256'hFFFFFEA525F4FFFF6867797F7EF3F354C1434646D1D5D4D45454D4D4D4D45554),
    .INIT_16(256'h54D4D4D4D623A45D7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFF7FFFFEA525737FFFFFFFFF7FFFEE6E42242A545455D5D454D5D5D5D5),
    .INIT_18(256'hCF4F4FCF4F4FCE4FD024A45D7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFF7BFB7B252472FFFEFEFFFFFFFF6D6E462C3155D554545450),
    .INIT_1A(256'hD5D55029A6A7A7A7A726A727A72424DE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFF7FFF26A425A4A4A4A5A5A5252525252525C35354D455),
    .INIT_1C(256'hD4D553D55454D0A62424A5A4A4A4A425A525A5DDFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFA7A3A4A4A42423A4A4A4A5A5A5A525C3),
    .INIT_1E(256'h9797182D3B3FD655463BBADFDFE56CEC6C6CEBEBEC5EDD463939FFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7939391D1897979798989898979797),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_001024_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n369,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_017,inst_doa_i1_016,inst_doa_i1_015,inst_doa_i1_014,inst_doa_i1_013,inst_doa_i1_012,inst_doa_i1_011,inst_doa_i1_010,inst_doa_i1_009}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h3FEFFFFFFFFFCA5F7EFFFFECB000E85FEFFFFF810025477AFFFFF838011336BF),
    .INITP_01(256'h00FF5FC7FFFFFCFFC1F07E7FFFFF87FC1FA239FFFFFE7FEDF25E9FFFFFC00261),
    .INITP_02(256'hFFFFFFFFB7FFFFFFFCFFDD4B7FFFFFFFE7FCE05FDFFFFFF9FFF1FFFF7FFFFFB8),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFF),
    .INIT_00(256'h000000000000002D57514644505455DCDEEEFFFFFFFFFFFEFFDCDD865553FFFF),
    .INIT_01(256'h5553FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFF154562102000200000000),
    .INIT_02(256'h090909090909090909090822434044464D5055DCE1EFFFFFFFFFFFFFFFDEDD85),
    .INIT_03(256'hFFFFFF935553FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF054541C0A070B),
    .INIT_04(256'h5850525555545454545454545454512A000956564B3C425754BEFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFF935553FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFF5659595553545555545554545554542600065650453E445455BEFFFF),
    .INIT_07(256'h4760716FE1E3EEFFFFFFFF955554FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFF5551431B1A1B1B1B1B1B1B1B1B1B192A38354746413E4046),
    .INIT_09(256'h3E3E3E3E3C4A5553DFDDEAFFFFFFFF955453FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFF5455420003010101010101010101002852523D3E),
    .INIT_0B(256'h554B3C3E3E3E3E3E3E495554E1DFECFFFFFFFF935251FFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55523E0C0D0B0B0B0B0B0B0B0B0B0B2E),
    .INIT_0D(256'h5555584A3E3B403E3E3E3E3E3E49555455555555555555C0FFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFEFF555255555555555555),
    .INIT_0F(256'h5454545454545648423E3E3E3E3E3E3E3E49555555555555555556BFFEFEFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF5854545454),
    .INIT_11(256'hD3D4D4D4D4D4D4D4D4D4D36E50505051515151515192D4D4D4D4D4D4D4D4D4EE),
    .INIT_12(256'hFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD4),
    .INIT_13(256'hFFFFFEFEFEFFFFFFFFFFFFFFFFFFFF78555556555555555556A9FFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFEFEFFFFFFFFFFFFFFFFFFFFFF78545555555455545455AAFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFEFEFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFDFBFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n412,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_008,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  // address_offset=2048;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hD1F3FFFFFD7FCC7FFFFFFFFF67FC06BFFFFFFF9E7FFF77FDFFFFF81FFEA13F9F),
    .INITP_01(256'hFFFFA7DFFFFFFEFFDDFFFAFFFFFFEFFE1FF3F7FFFFF3FFEFFFBF3FFFFF380197),
    .INITP_02(256'hFFFFFDFFFFFFFFFFFFFFEDFFFFFFFFFFFFFF9F7FDFFFFFFE0009F801FFFFFF67),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFBFFFFFF),
    .INIT_00(256'h0C0C0C0C0C0C0C17A429555437A5A56EEFF77FFFFFFFFF7FFF6EEEC0A4A4FFFF),
    .INIT_01(256'hA4A4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF72525168C8C8A8B0C0C0C),
    .INIT_02(256'h8E0E0E0E0E0E0E0E0E0E8E179FA6D151B928A9EF6E76FFFFFFFFFFFFFF6FEE40),
    .INIT_03(256'hFFFFFFC7A4A4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF7A525968E0E0E),
    .INIT_04(256'h25A625A4A525A52525A52525A525A5970C0E25A5B9C542A7255CFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFC7A4A4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFF7FFFA5A4A323A4A3A3A3A3A3A3A3A3A323188C8E2425BA43C027A5DDFFFF),
    .INIT_07(256'hBBB934B4F0F0F6FFFFFFFFC7A4A4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFF2525A0949514141414141414141413171C1FBABCC14443BC),
    .INIT_09(256'hC3C3C3C3C4B4A4256EEE75FFFFFFFFC7A4A5FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFA5249C0C0C8B8B8B8B8B8B8B8B8B8C9825A843C3),
    .INIT_0B(256'hA8AC43C3C3C3C3C3C3B4A425EDEEF47F7FFFFEC7A526FFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA5259F8F908F8F8F8F8F8F8F8F8F909B),
    .INIT_0D(256'hA4A4A3B5C4C4C4C3C3C3C3C344B425A525A4A4A4A4A4A55DFF7FFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7E7FFFA5A4A4A4A4A4A4A4A4),
    .INIT_0F(256'h25252525252524B543C3C3C3C3C3C3C344B325A4A4A4A4A4A4A4A5DD7F7FFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEA5A4252525),
    .INIT_11(256'h68E8E8E8E8E8E8E8E8E868372B2BAB2A2A2A2A2AAA4968E8E8E8E8E8E8E8E8F6),
    .INIT_12(256'hFFFF7EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8),
    .INIT_13(256'hFFFF7EFFFFFFFFFFFFFFFFFFFFFFFFB8A424242525252525A551FFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFF7F7FFFFFFFFFFFFFFFFFFFFF7F382424A5A4A5A4A5A524D27F7F),
    .INIT_16(256'h7E7F7FFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFF7EFEFF7FFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFF7FFEFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFD7F7FFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_002048_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n455,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_017,inst_doa_i2_016,inst_doa_i2_015,inst_doa_i2_014,inst_doa_i2_013,inst_doa_i2_012,inst_doa_i2_011,inst_doa_i2_010,inst_doa_i2_009}));
  // address_offset=3072;data_offset=0;depth=528;width=9;num_section=1;width_per_section=9;section_size=24;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'h000000000000000000000000000000000000000000000000000000000000FFFF),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_3600x24_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({open_n498,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_008,inst_doa_i3_007,inst_doa_i3_006,inst_doa_i3_005,inst_doa_i3_004,inst_doa_i3_003,inst_doa_i3_002,inst_doa_i3_001,inst_doa_i3_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i1_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_1  (
    .i0(inst_doa_i2_010),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b10/B0_0 ),
    .i1(\inst_doa_mux_b10/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_0  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i1_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_1  (
    .i0(inst_doa_i2_011),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b11/B0_0 ),
    .i1(\inst_doa_mux_b11/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_0  (
    .i0(inst_doa_i0_012),
    .i1(inst_doa_i1_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_1  (
    .i0(inst_doa_i2_012),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b12/B0_0 ),
    .i1(\inst_doa_mux_b12/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[12]));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_0  (
    .i0(inst_doa_i0_013),
    .i1(inst_doa_i1_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_1  (
    .i0(inst_doa_i2_013),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b13/B0_0 ),
    .i1(\inst_doa_mux_b13/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[13]));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_0  (
    .i0(inst_doa_i0_014),
    .i1(inst_doa_i1_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_1  (
    .i0(inst_doa_i2_014),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b14/B0_0 ),
    .i1(\inst_doa_mux_b14/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[14]));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_0  (
    .i0(inst_doa_i0_015),
    .i1(inst_doa_i1_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_1  (
    .i0(inst_doa_i2_015),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b15/B0_0 ),
    .i1(\inst_doa_mux_b15/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[15]));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_0  (
    .i0(inst_doa_i0_016),
    .i1(inst_doa_i1_016),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_0 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_1  (
    .i0(inst_doa_i2_016),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_1 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b16/B0_0 ),
    .i1(\inst_doa_mux_b16/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[16]));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_0  (
    .i0(inst_doa_i0_017),
    .i1(inst_doa_i1_017),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_0 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_1  (
    .i0(inst_doa_i2_017),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_1 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b17/B0_0 ),
    .i1(\inst_doa_mux_b17/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[17]));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_0  (
    .i0(inst_doa_i0_018),
    .i1(inst_doa_i0_018),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_0 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_1  (
    .i0(inst_doa_i0_018),
    .i1(inst_doa_i0_018),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_1 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b18/B0_0 ),
    .i1(\inst_doa_mux_b18/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[18]));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_0  (
    .i0(inst_doa_i0_019),
    .i1(inst_doa_i0_019),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_0 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_1  (
    .i0(inst_doa_i0_019),
    .i1(inst_doa_i0_019),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b19/B0_1 ));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b19/B0_0 ),
    .i1(\inst_doa_mux_b19/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[19]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_0  (
    .i0(inst_doa_i0_020),
    .i1(inst_doa_i0_020),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_0 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_1  (
    .i0(inst_doa_i0_020),
    .i1(inst_doa_i0_020),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b20/B0_1 ));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b20/B0_0 ),
    .i1(\inst_doa_mux_b20/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[20]));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_0  (
    .i0(inst_doa_i0_021),
    .i1(inst_doa_i0_021),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_0 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_1  (
    .i0(inst_doa_i0_021),
    .i1(inst_doa_i0_021),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b21/B0_1 ));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b21/B0_0 ),
    .i1(\inst_doa_mux_b21/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[21]));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_0  (
    .i0(inst_doa_i0_022),
    .i1(inst_doa_i0_022),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_0 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_1  (
    .i0(inst_doa_i0_022),
    .i1(inst_doa_i0_022),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b22/B0_1 ));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b22/B0_0 ),
    .i1(\inst_doa_mux_b22/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[22]));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_0  (
    .i0(inst_doa_i0_023),
    .i1(inst_doa_i0_023),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_0 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_1  (
    .i0(inst_doa_i0_023),
    .i1(inst_doa_i0_023),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b23/B0_1 ));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b23/B0_0 ),
    .i1(\inst_doa_mux_b23/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[23]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i1_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_1  (
    .i0(inst_doa_i2_009),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b9/B0_0 ),
    .i1(\inst_doa_mux_b9/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[9]));

endmodule 

