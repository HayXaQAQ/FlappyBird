// Verilog netlist created by TD v4.6.18154
// Wed Nov 11 23:52:47 2020

`timescale 1ns / 1ps
module ggbutton  // al_ip/ygyhu.v(14)
  (
  addra,
  addrb,
  clka,
  clkb,
  rsta,
  rstb,
  doa,
  dob
  );

  input [12:0] addra;  // al_ip/ygyhu.v(21)
  input [12:0] addrb;  // al_ip/ygyhu.v(22)
  input clka;  // al_ip/ygyhu.v(23)
  input clkb;  // al_ip/ygyhu.v(24)
  input rsta;  // al_ip/ygyhu.v(25)
  input rstb;  // al_ip/ygyhu.v(26)
  output [7:0] doa;  // al_ip/ygyhu.v(18)
  output [7:0] dob;  // al_ip/ygyhu.v(19)

  wire [0:0] addra_piped;
  wire [0:0] addrb_piped;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_dob_i0_000;
  wire inst_dob_i0_001;
  wire inst_dob_i0_002;
  wire inst_dob_i0_003;
  wire inst_dob_i0_004;
  wire inst_dob_i0_005;
  wire inst_dob_i0_006;
  wire inst_dob_i0_007;
  wire inst_dob_i1_000;
  wire inst_dob_i1_001;
  wire inst_dob_i1_002;
  wire inst_dob_i1_003;
  wire inst_dob_i1_004;
  wire inst_dob_i1_005;
  wire inst_dob_i1_006;
  wire inst_dob_i1_007;

  reg_sr_as_w1 addra_pipe (
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped));
  reg_sr_as_w1 addrb_pipe (
    .clk(clkb),
    .d(addrb[12]),
    .en(1'b1),
    .reset(rstb),
    .set(1'b0),
    .q(addrb_piped));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CSAMUX("INV"),
    .CSBMUX("INV"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h202020202020202020202020202020202121212121201F1F1901010102040603),
    .INIT_01(256'h2020202020202020202020202020202020202020202020202020202020202020),
    .INIT_02(256'h201F1E1F20211F1F202020202020202020202020202020202020202020202020),
    .INIT_03(256'h010101010101010101010101020202010101000003000003020201012021201F),
    .INIT_04(256'h0101010101010101010101010101010101010101010101010101010101010101),
    .INIT_05(256'h0202020101000000000000010101010101010101010101010101010101010101),
    .INIT_06(256'h0404040404040404050504040404040403030201010202050000000000000101),
    .INIT_07(256'h0404040404040404040404040404040404040404040404040404040404040404),
    .INIT_08(256'h0403030303040404040404040404040404040404040404040404040404040404),
    .INIT_09(256'h0E0E0E0F0F0F0E0F10100F0F0E0D0A0702000102000000020203040404050404),
    .INIT_0A(256'h0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E),
    .INIT_0B(256'h0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E),
    .INIT_0C(256'h2828272729292828292A322D09030501000001040A0D0E0E0E0F0E0E0E0E0E0E),
    .INIT_0D(256'h2828282828282828282828282828282828282828282828282828282828282828),
    .INIT_0E(256'h2828282828282828282828282828282828282828282828282828282828282828),
    .INIT_0F(256'h3536353534313A360A0402000101030A1D242726272828272827272727282828),
    .INIT_10(256'h3435343534353435343534353435343534353435343534353435343435353334),
    .INIT_11(256'h3435343534353435343534353435343534353435343534353435343534353435),
    .INIT_12(256'h3A3434310A0202000101040D2730333332353435343534353435343534353435),
    .INIT_13(256'h3636363636363636363636363636363636363636363636363736353537373636),
    .INIT_14(256'h3636363636363636363636363636363636363636363636363636363636363636),
    .INIT_15(256'h0A0000030101050E283136363436373636363636363636363636363636363636),
    .INIT_16(256'h3636363636363636363636363636363636363637383736363737363633373732),
    .INIT_17(256'h3636363636363636363636363636363636363636363636363636363636363636),
    .INIT_18(256'h0102040F29333937353638373636363636363737363636363636363636363636),
    .INIT_19(256'h3737373737373737373737373737373839383636373736363637383608000001),
    .INIT_1A(256'h3737373737373737373737373737373737373737373737373737373737373737),
    .INIT_1B(256'h2736363638363837373737373737373737373737373737373737373737373737),
    .INIT_1C(256'h3737373737373737373737383939363637373636363739360800000102020310),
    .INIT_1D(256'h3737373737373737373737373737373737373737373737373737373737373737),
    .INIT_1E(256'h3837383737373737373737373737373737373737373737373737373737373737),
    .INIT_1F(256'h3737373737373737383836373737363636373836070001020202031027363636),
    .INIT_20(256'h3737373737373737373737373737373737373737373737373737373737373737),
    .INIT_21(256'h3737363636373737373737373737373737373737373737373737373737373737),
    .INIT_22(256'h3637363737373737373736363636383607000102020203102735363637363837),
    .INIT_23(256'h3637363736373637363736373637363736373637363736373637363736373637),
    .INIT_24(256'h3636363636373637363736373637363736373637363736373637363736373637),
    .INIT_25(256'h3737383837373636363637360700010202020310273536363736383737373636),
    .INIT_26(256'h3737373737373737373737373737373737373737373737373737373737373737),
    .INIT_27(256'h3737373737373737373737373737373737373737373737373737373737373737),
    .INIT_28(256'h3737373736363735070001020202031027353636373638373737373737373737),
    .INIT_29(256'h3737373737373737373737373737373737373737373737373737373736373838),
    .INIT_2A(256'h3737373737373737373737373737373737373737373737373737373737373737),
    .INIT_2B(256'h3636363406000001020203102736363638363837373737373637363737373737),
    .INIT_2C(256'h3636363636363636363636363636363636363636363636363636373736373737),
    .INIT_2D(256'h3636363636363636363636363636363636363636363636363636363636363636),
    .INIT_2E(256'h0600000001020310273535353736373736363636363636363636363636363636),
    .INIT_2F(256'h3536363736363636363736363535353636363737353636373636373736363634),
    .INIT_30(256'h3736363637373636363637373737373636363737373737373636363636363535),
    .INIT_31(256'h0102031027353536373537363636363636373737373735353636363636363637),
    .INIT_32(256'h36393937383A39343235343537393D3939363637353638373737363407000000),
    .INIT_33(256'h393C3C39373638383A38373637393C413D3C3B39363435363636373532343937),
    .INIT_34(256'h263335373735373937373839393A3C3B3A3834343838383A3834373939383736),
    .INIT_35(256'h3E42444343474344454547413E39363734343838383836350701000002020410),
    .INIT_36(256'h3836373737383739414D53514D48413D3937393D4342403B343539383737393B),
    .INIT_37(256'h3835363637393C40424445474646424246443E3A363435393A393A415150493F),
    .INIT_38(256'h5C5F5C5C5B58574E403B38373434383838383635070100000202041026333437),
    .INIT_39(256'h35393838475F67615B564F494444484D595750463D393A39393B414C5356595D),
    .INIT_3A(256'h3B444E55585A5B5D5C5D5A5859554A403737353739383D4E656258483D373535),
    .INIT_3B(256'h69655E52413B38363434383838383635080100000202040F2733353738343435),
    .INIT_3C(256'h4258626062605F5D5B5A5D6167665E4F423938393D47545E6161626261666567),
    .INIT_3D(256'h64605E5F64656765635E52433839363639373D5765645D514339353536393737),
    .INIT_3E(256'h403A36363435373738383634080100000202040F283435373733383C4E555F64),
    .INIT_3F(256'h575A5C5E5D5D5F62656961514336333A4858646057524F4A4C53555F67655C4D),
    .INIT_40(256'h54586166625C4E3F373936363937405B60636157493B35333436353539434C4F),
    .INIT_41(256'h353637373837363408010000020204102735373736343E4A5D5F5E59514B4747),
    .INIT_42(256'h4443464B5D655F514335334054616454433D3A37393D415161645A4A3F393535),
    .INIT_43(256'h61584B3B36373535383B485F6364635D4F413835333538383737383D3F404344),
    .INIT_44(256'h3837363408010000020204102735373736374859645D50433B38393A3F445665),
    .INIT_45(256'h58645F53443938495D615C4A39353536363738485E645D4C403A353635363737),
    .INIT_46(256'h37353536383F526462605F5F594D423B3636383A3936333636383A3B3B3B3F42),
    .INIT_47(256'h080000000202041027343536363A50636457453A36373B3C38394D6161584A3B),
    .INIT_48(256'h463A3C4E6561584739343638393734445B655E4C423B36363536383738373634),
    .INIT_49(256'h374358675A58585E5F574A423A38373739393636424446484846484C58656454),
    .INIT_4A(256'h0202041027323336383E55686254413735373C3C3935475E60594D3E39363635),
    .INIT_4B(256'h61625E4D3D38393A3836353F55666155453C3537363638383837353308000001),
    .INIT_4C(256'h574C47556260554A3F3935373836383F57595B5D5E5E5D5C60636056473B3E4E),
    .INIT_4D(256'h25343534374258676157473A36383D3C393B435C665C4E4237363A36364B6264),
    .INIT_4E(256'h443E3B3A3836353D52646053453C353836363837373735330800000102020410),
    .INIT_4F(256'h5B635D53463D36343534383F5456585A5D5D5E5E5F646459493D3C4662625E51),
    .INIT_50(256'h363C5062645C4F4038373A3A393A435B675E50433B3735343D546461584B424A),
    .INIT_51(256'h383734394D636356473D36363636383737373534080000010202041027343536),
    .INIT_52(256'h504338333433363B4143424444454545525E625B4C403B3E595E625B4E443E39),
    .INIT_53(256'h6360574B3F39383736373E56666054453B373336475D65615C51474A5761615D),
    .INIT_54(256'h4860645A4A3E3736363638383737353408000001020204102A35363937374657),
    .INIT_55(256'h333335383A3A3736343535354356625D5042393947546164594D44403C3A3537),
    .INIT_56(256'h4B433D3A3636394E636358473937343A4F6065635F5D5B5A5C616363584C3D36),
    .INIT_57(256'h4C3F3737353638373736353308000101020204102835383937343D485D605E56),
    .INIT_58(256'h3E3E3B3A3939393940576663554338353945565F605B565248463F3D485C625C),
    .INIT_59(256'h3F3B394C61655B49393635405663625E5B5F6361606365676156463A35363A3D),
    .INIT_5A(256'h3537383737363533080001010202040F26363636353538384E5861625C534B45),
    .INIT_5B(256'h42403F404255646458473A36373B43505B6163615A58504B525F635F50413837),
    .INIT_5C(256'h63655C4A3D3638495F655C504E505256595E6367665E4E3F383B434A48464543),
    .INIT_5D(256'h37363433080001010202040F24353635363738333B47576063625D574F4C4652),
    .INIT_5E(256'h4C5961625B4C3D3839393A4049535A5E61615E5C5E6365615241383635363837),
    .INIT_5F(256'h403941566361534341414244464A545D636157493F4450595857565453525150),
    .INIT_60(256'h07000102020204102634353738373735363B444D575E62615D5C565D66665E4E),
    .INIT_61(256'h5E4D3D3738383838393E4A545E5F616263646361544337363636373736363533),
    .INIT_62(256'h63594B3D393B3B3A363742525E625F53494C5862606060606160605F5D626363),
    .INIT_63(256'h0202041028333538393638393939383B4350595C6164616468655E4F3F3B4D61),
    .INIT_64(256'h3737373637373A3B474E565D6569635A4C413735363433343636363507010101),
    .INIT_65(256'h37383A39383A3C3E555E645E51494B52585757595A5D5F61616468675A463B37),
    .INIT_66(256'h273536363737383738383738393E444755595F63676456473A44576562514039),
    .INIT_67(256'h36373839393E444B545A5751433C363637363536353739360700000101020310),
    .INIT_68(256'h37383A3C454F59574B403C3C403F414245484C4D525558584E40383737363636),
    .INIT_69(256'h37363737383736363537393B3A434F575C594A3D373D4B565347393535373838),
    .INIT_6A(256'h3536373A3F43423E3A3734363937363837383A36080000010102031027353536),
    .INIT_6B(256'h383D43423C3836373737363635383A3C3F4042433E3735363636373636373637),
    .INIT_6C(256'h373738373636363732373D4144453D3534373E44423933333436373736363639),
    .INIT_6D(256'h35373633363534373837363838393936080101020102030F2735363637363837),
    .INIT_6E(256'h3537373A38383636343436373737393937343437363736373736363636363635),
    .INIT_6F(256'h3738383837383737373836353636373938353335343637363636363636373736),
    .INIT_70(256'h353536373736353736373735070002030102030F273535363735373736363738),
    .INIT_71(256'h38373735363737383838393A3837363836363638373737373838363535373533),
    .INIT_72(256'h3637393838383737383737373736353735363638373737373737383738383737),
    .INIT_73(256'h3737363737363735070103040102030F27353636373638373738383837363637),
    .INIT_74(256'h3737373739383939383735363636373738383837363737373637373734353737),
    .INIT_75(256'h3838383938383738373737373536363838383838383837373837383738373637),
    .INIT_76(256'h36363735080103040102030F2736363638373837373838373637373737383839),
    .INIT_77(256'h3737363637363534353636363738383838383939383737373536373738383637),
    .INIT_78(256'h363736363537363636363637373837373837363536363A3A3937373737363636),
    .INIT_79(256'h08010202010203102736363638373838373737373738393A3A39363535353638),
    .INIT_7A(256'h3839373636363636373738393739393837373739363738373838353536363735),
    .INIT_7B(256'h3637383737363535373737363537393737363637363635363636363637383738),
    .INIT_7C(256'h0102031027363636383738373737373736373737373736383837373737373635),
    .INIT_7D(256'h3535353536363637373737373736363637373838373736363738373207000001),
    .INIT_7E(256'h3736373737373737373636363636363637393838383838383939393938383737),
    .INIT_7F(256'h27333633363837353636363636363637393937373637393A3A3937373737393A),
    .MODE("DP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_5000x8_sub_000000_000 (
    .addra(addra[11:1]),
    .addrb(addrb[11:1]),
    .bytea(addra[0]),
    .byteb(addrb[0]),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12]),
    .csb(addrb[12]),
    .dia({open_n49,open_n50,open_n51,open_n52,open_n53,open_n54,open_n55,open_n56,8'b00000000}),
    .dib({open_n57,open_n58,open_n59,open_n60,open_n61,open_n62,open_n63,open_n64,8'b00000000}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({open_n69,open_n70,open_n71,open_n72,open_n73,open_n74,open_n75,open_n76,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}),
    .dob({open_n77,open_n78,open_n79,open_n80,open_n81,open_n82,open_n83,open_n84,inst_dob_i0_007,inst_dob_i0_006,inst_dob_i0_005,inst_dob_i0_004,inst_dob_i0_003,inst_dob_i0_002,inst_dob_i0_001,inst_dob_i0_000}));
  // address_offset=4096;data_offset=0;depth=904;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h373737383838373737373636373839393838373739383633080102030202030F),
    .INIT_01(256'h3838383837373737373736373839393939393939393939393939383837373636),
    .INIT_02(256'h353836353736363636373738393938383738393A3A39383838383A3A38383838),
    .INIT_03(256'h363636363535353536373738383838393A3A3A37090001020202030F28333734),
    .INIT_04(256'h3636363635353535363636373737373737373737373736363737373737373737),
    .INIT_05(256'h3636363636363637373736363636373838373636363638383636363637373636),
    .INIT_06(256'h3636363636373838383838393C383437090604010202030F2733383535363535),
    .INIT_07(256'h3636363636363636363636373636363636363637383939383838383837373636),
    .INIT_08(256'h3737373737373635353636373736363636363737373838383737373737373736),
    .INIT_09(256'h343435353535353635363836090302020102030F273338363636363737373737),
    .INIT_0A(256'h3332333333333333333332333333333436363636363535353535353535353534),
    .INIT_0B(256'h3433333232323333333332323233333435353535353535353535353535353434),
    .INIT_0C(256'h262526262B2F342F070104060202030E26323534353534363535353535353535),
    .INIT_0D(256'h2525252424252524252525252727272727262626262626262627262625252727),
    .INIT_0E(256'h2425252525252425242525262627272726272727272727272726262625252525),
    .INIT_0F(256'h0D0A0906000502020202030B1C23262528282729272626262626262626262525),
    .INIT_10(256'h10100F1010111111100F0F0F0F0F0F0F0F1010111112121210111312100F0F0E),
    .INIT_11(256'h1010101010111110100F0F100F10101010111010100F0F0F1011101111111111),
    .INIT_12(256'h01020203020202060A0F0E0E10111010101010100F1010111112111110101010),
    .INIT_13(256'h0404040403020202020202020202030304050504040406050302010202030401),
    .INIT_14(256'h0404040403020303030303030302020202020303030404040504050404040304),
    .INIT_15(256'h0201020202020202030403030403030303030304040504040404040404040404),
    .INIT_16(256'h0808080707070707070808080808080808080808080707070708010001020000),
    .INIT_17(256'h0808080808080808080808080808080808080808080808080808080808080808),
    .INIT_18(256'h0707080808080808080808080808080808080808080808080808080808080808),
    .INIT_19(256'h19191919191919191919191919191919191919191A1802020000000008080808),
    .INIT_1A(256'h1919191919191919191919191919191919191919191919191919191919191919),
    .INIT_1B(256'h1919191919191919191919191919191919191919191919191919191919191919),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000001919191919191919),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_5000x8_sub_004096_000 (
    .addra(addra[11:1]),
    .addrb(addrb[11:1]),
    .bytea(addra[0]),
    .byteb(addrb[0]),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[12]),
    .csb(addrb[12]),
    .dia({open_n87,open_n88,open_n89,open_n90,open_n91,open_n92,open_n93,open_n94,8'b00000000}),
    .dib({open_n95,open_n96,open_n97,open_n98,open_n99,open_n100,open_n101,open_n102,8'b00000000}),
    .rsta(rsta),
    .rstb(rstb),
    .doa({open_n107,open_n108,open_n109,open_n110,open_n111,open_n112,open_n113,open_n114,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}),
    .dob({open_n115,open_n116,open_n117,open_n118,open_n119,open_n120,open_n121,open_n122,inst_dob_i1_007,inst_dob_i1_006,inst_dob_i1_005,inst_dob_i1_004,inst_dob_i1_003,inst_dob_i1_002,inst_dob_i1_001,inst_dob_i1_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped),
    .o(doa[7]));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_0_0  (
    .i0(inst_dob_i0_000),
    .i1(inst_dob_i1_000),
    .sel(addrb_piped),
    .o(dob[0]));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_0_0  (
    .i0(inst_dob_i0_001),
    .i1(inst_dob_i1_001),
    .sel(addrb_piped),
    .o(dob[1]));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_0_0  (
    .i0(inst_dob_i0_002),
    .i1(inst_dob_i1_002),
    .sel(addrb_piped),
    .o(dob[2]));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_0_0  (
    .i0(inst_dob_i0_003),
    .i1(inst_dob_i1_003),
    .sel(addrb_piped),
    .o(dob[3]));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_0_0  (
    .i0(inst_dob_i0_004),
    .i1(inst_dob_i1_004),
    .sel(addrb_piped),
    .o(dob[4]));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_0_0  (
    .i0(inst_dob_i0_005),
    .i1(inst_dob_i1_005),
    .sel(addrb_piped),
    .o(dob[5]));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_0_0  (
    .i0(inst_dob_i0_006),
    .i1(inst_dob_i1_006),
    .sel(addrb_piped),
    .o(dob[6]));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_0_0  (
    .i0(inst_dob_i0_007),
    .i1(inst_dob_i1_007),
    .sel(addrb_piped),
    .o(dob[7]));

endmodule 

