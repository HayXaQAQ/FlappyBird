// Verilog netlist created by TD v4.6.18154
// Sat Nov 14 16:30:10 2020

`timescale 1ns / 1ps
module grass  // al_ip/star.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [12:0] addra;  // al_ip/star.v(18)
  input clka;  // al_ip/star.v(19)
  input rsta;  // al_ip/star.v(20)
  output [7:0] doa;  // al_ip/star.v(16)

  wire [0:0] addra_piped;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;

  reg_sr_as_w1 addra_pipe (
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSAMUX("INV"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_01(256'hFAF5FAFAF6F4B880808080808080808080808080808080808080808080808080),
    .INIT_02(256'h80808080808BB2F2ECE8E9EFF1F9F3B9898080808080808080808080B2FDFBFB),
    .INIT_03(256'hACA7AA8080808080808080808080808080808080808080808080808080808080),
    .INIT_04(256'hF4F7E4B180808080808080808080808080808080808080808080808789ACA5A9),
    .INIT_05(256'h86AFE8ECE0E5DFE0E7EFF2DFAE80808080808080808080AEEDF8F5F2E7E4EEF3),
    .INIT_06(256'h8080808080808080808080808A80808080808080808080808080808080808080),
    .INIT_07(256'h80808080808080808080808080808080808080808080AA91BBE8E2EFF3EBE8B2),
    .INIT_08(256'hDDDAD3D6DFE5EDECEEA68080808080808080A6E7F3EAE6DDE2DFE7EFEEEDEEA7),
    .INIT_09(256'h80808080808081A4A3B0B38680808080808080808080808080808080A6E9F6E5),
    .INIT_0A(256'h8080808080808080808080808080849894D5CEA0E6ECE2DCE2EDF1E4A98B8080),
    .INIT_0B(256'hD6DDE7E3E7F2AB80808080808080AFF2EBE8DCDDDCDADFE9EBE6EB8080808080),
    .INIT_0C(256'h81ADAAD7EEE7E3B08E808080808080808080808080808080B2F7E6E0E0D2D4DB),
    .INIT_0D(256'h8080808080808080818983A1A1ABACC2E1D9DEDCE0E6E2E7E7A3888080808080),
    .INIT_0E(256'hEBEDA4808080808080A8E5E9E4E5DFDDD9DCDDE5E8E6E2808080808080808080),
    .INIT_0F(256'hEAE7DBE2A4898080808080808080808080808088ACE6E4DBD9D2D9D8CFD5DFE4),
    .INIT_10(256'h8080808B8B9B979F999C95DADBDCDCDFE1E1E4E5F0AB868080808080ABC0D5CF),
    .INIT_11(256'h808080808080B4ECEDDED9DEDEE0DEDDE1E2CB80808080808080808080808080),
    .INIT_12(256'hAD8D8080808080808080808080808080B3EFE2DCD2D8D8D2D7D9D5DEEAE9B380),
    .INIT_13(256'h95969497A191CFD9D6DBD8DCDFE0E4DFDCBB80808080809CACD5D8DAD1D8D2D7),
    .INIT_14(256'h8080A2E9E2DEDDD8DADFDDDEE5EAB9A58080808080808080808080808080809B),
    .INIT_15(256'h808080808080808080808080ACE5E3E0D7D7D5D4DEDECFD6DEBB808080808080),
    .INIT_16(256'h8A82DFE6DBD9DADBDDE0DEDFE6E08080808080A6D4D8D8CCD4D6D8CACCA68080),
    .INIT_17(256'hD4DFDFD5DDDDDBE1ECEEA7B5928080808080808080808080808D979498959598),
    .INIT_18(256'h808080808080808089B0EFE1DBD1DCDDD7D7D5D8E7E280808080808080808DB3),
    .INIT_19(256'hE1E1DAD6DADDDED8DEB5979980808082B9DCD4D1D2DAD8D4D0DAAA8080808080),
    .INIT_1A(256'hE0DCDDB0AFDF7E94B5808080808080808080807E8A98928E9490949D97B5F2E2),
    .INIT_1B(256'h80808080808CABE9E2D7DDE1E4DCD9E2AB80828080808080808080A6B1D4DCE1),
    .INIT_1C(256'hDBD0D3DEB98FDA8980808080B1EAD4DADBD4D9D7D3D2A1808080808080808080),
    .INIT_1D(256'h80808FA789808080808080808080978F9891908E9296968B89E7E9E2DEDBD7DC),
    .INIT_1E(256'h8085B3ECE6E5E9E7E4DEB6A7808080808A8080808080808080B4E4E9E2DCAC8F),
    .INIT_1F(256'h7890CC808080808086B1DFDAD9D9D9D7D1D7AB80808080808080808080808080),
    .INIT_20(256'h988B808080808080809D9F9B9F96918F90959A86ADECE4E1E1E2D9DADBD7E8D3),
    .INIT_21(256'hEFE6EEE5E4AC8B8080808980B5988080808080808080E5EEE2AD808080808098),
    .INIT_22(256'h808080808AABDFD4DBCEDACECBCEAA808080808080808080A397838080808FAF),
    .INIT_23(256'h80808080808089857C84959496999C9388E0E9DFDBE2E0E0E0DDE2948BA19580),
    .INIT_24(256'hAE808080808080808EA696848A8080808A8090C1A98080808080809095878080),
    .INIT_25(256'h80A2E1D0CDCDC9C9B2A68980808080808080808080809992828080DCE4EFA6AC),
    .INIT_26(256'h9380A78B80868382869C8B8080A8F2E3E8E7E4E6E3E6C498A29E8B8080808080),
    .INIT_27(256'h80808080979E98877E808080808098779A808080808093949680808080808080),
    .INIT_28(256'hBFA6BFAC8D8080808080808080808080809AA097868992899980808080808080),
    .INIT_29(256'h9D9885847C8B88808088A8F0EDEDEBEAEAE684899B93908080808080808DA7DF),
    .INIT_2A(256'h828F969B8C878080809AA68E958680808080809995878080808080929D899399),
    .INIT_2B(256'h808080808080808080808080808E95969C9B95848B928A808080808080808080),
    .INIT_2C(256'h7F8C808080808CAEEEF2E9E3F0D58E9E949E8D8080808080808088A9A0C1BF88),
    .INIT_2D(256'h928B808080939D989B8982808080889B929B8D808080808B9D8480979A939696),
    .INIT_2E(256'h80808080808080808084869B99929D97959A8982808A8080808080808A88998E),
    .INIT_2F(256'h808080ADEDF0F0EEEA958E959B8680808080808080808091AA97808080808080),
    .INIT_30(256'h80919C93979D898080838E9998988D8080808B9A95A08A778A96929696998A80),
    .INIT_31(256'h808080808080879B9797929694949C888C818980808080808A90999391968F80),
    .INIT_32(256'h9BA5ACA4D78384969B8A80808080808080808A9C998F80808080808080808080),
    .INIT_33(256'h9694A18C847C8995919790808080889698979D837C87969393979B8780808088),
    .INIT_34(256'h8080808B969291929293939594878B8A8080808080808A93918E9B9291909B8F),
    .INIT_35(256'h808FA096978D80808080808080989C9299898080808080808080808080808080),
    .INIT_36(256'h8689989196968580808089999790979B8C888595959896968091808080868086),
    .INIT_37(256'h9C95909293929091928E988B8289808080808A9992919389828D929091959285),
    .INIT_38(256'h978C808080808080918C939C8B8080808080879D80808080808080808080808A),
    .INIT_39(256'h919A9A8080807C9696949499997C899B9693979A9B9E90808080808080929797),
    .INIT_3A(256'h9795929293939B958A8D808A808089A09195949C8888998E8F92959B7D89979A),
    .INIT_3B(256'h8080808A9597979A8D8080808580AF8080808080808080808080808087969997),
    .INIT_3C(256'hA199A19A9494948F91998A839C97938E9594999280808080868D9F9799868080),
    .INIT_3D(256'h9393979293998F8180808A8C97949799887B82928B8E96988A889C95968F968B),
    .INIT_3E(256'h988F958280808080809BBE808080808080808080808080808D99978C95959293),
    .INIT_3F(256'h918F92918E99838584979394919698A0928080807A899B91988080808080838C),
    .INIT_40(256'h9990968B8A8080929C8E9497978A7A98978F9697807C7E94918E9B86898B9D94),
    .INIT_41(256'h8080808089C08080808080808080808080808080808594958E91919494949693),
    .INIT_42(256'h91909B8880859592919191968C8480888E99939E97858080808080989293988E),
    .INIT_43(256'h93808085859495909096858C969791908A8B9D94919397858A919D9591909293),
    .INIT_44(256'h95B68080808080808080808080808080808F968C8F9191949397949592978F9B),
    .INIT_45(256'h89839991958E95948E888080879E939598888080808A9E9F999A9B8A80808080),
    .INIT_46(256'h849995919590847988938E938983969491949A8C81919B91919493919493A09D),
    .INIT_47(256'h808080808080808080808080808081959192929492948F948B9593949C8E8790),
    .INIT_48(256'h92959090858680808B949A9699878080808A9D92939A907F81808095AA908080),
    .INIT_49(256'h8C939B88849792918884989590909A857C869891919193979697818589818196),
    .INIT_4A(256'h808080808080808080808A979191919592958D9397949390949E938A8B94948E),
    .INIT_4B(256'h9B89809485939595978F808080869696939C8F8781908D9DA18E808080808080),
    .INIT_4C(256'h8A82969789849E928F9390948C968F9190939298959782899C87809D96938F91),
    .INIT_4D(256'h808080808080919B938894909293949292939494969898917E89938F8B909B99),
    .INIT_4E(256'h899A93919C8080808698978D959A94898993A1939C8B80808080808080808083),
    .INIT_4F(256'h8F8793958F9392948E948F90918E95938F847B8295837F8095948F90978DA48B),
    .INIT_50(256'h80807B8E979196939192939292939594959697978D8394929091979B8582819B),
    .INIT_51(256'h94808080909796938DA09B96888D9799998A8080808080808080808080969980),
    .INIT_52(256'h9193949391939392988F8F9A9184869B999B7C88999294989888817B89958D94),
    .INIT_53(256'h93959493919191908D9094949294989A827D818A8D8D92979D7F83A18C8C9E90),
    .INIT_54(256'h818E9294907A85A8939D9097978A8080808080808080808080A19A98947D8F8B),
    .INIT_55(256'h919195939191928D968E8296949387888F919793909D927585969090988B8081),
    .INIT_56(256'h9192918E8B8E9493919295989B7E989491908F9092827C90B4949D8F9393938E),
    .INIT_57(256'h938A99818A909394988B80808080808080808080809D9893968C8F7C85949194),
    .INIT_58(256'h959793919A838B99979494838594969596979C7E88938B949A89A8919D98958E),
    .INIT_59(256'h8F90929492939597999394908D939293969C8A9CBB89A0979693928D93929593),
    .INIT_5A(256'h96908E96988C8080808080808080808085939B9295949D878294919492929390),
    .INIT_5B(256'h8D7E8C9994979A8083978B95909889788094929098868E89968D92979686838E),
    .INIT_5C(256'h9293959596988E9192908F8F8E9D8C87B2989392949294909492949297928796),
    .INIT_5D(256'h988D8080808080808080808080968D908C8F9783849192939292939393919090),
    .INIT_5E(256'h969495837F9C9794939C859198888D96998C7E8899949296A2878B9C94909194),
    .INIT_5F(256'h8E9491949890939196929A8A9E9698949191949392909293969694968F7E7E86),
    .INIT_60(256'h8080808080808080848997988F8E9297838992919091939595938F8E92939191),
    .INIT_61(256'h7D829794928E867F989292939884869C989094998A7C7F9491918E93988F8080),
    .INIT_62(256'h948B9492939896868A899C9293939594919193969297919A8DA78C8597969C8A),
    .INIT_63(256'h80808080808A9796919290928284969393929393949592929593918F9193988F),
    .INIT_64(256'h93939595939292929081979594938F9A8884999391918F949C8A808080808080),
    .INIT_65(256'h939A947F7D829996959494949393959593949494888A9583829DA0857D8B9696),
    .INIT_66(256'h8090999595918B91977A83979298949595959494959492929291929292919293),
    .INIT_67(256'h93939392948994939495969981819493939190939B8D80808080808080808080),
    .INIT_68(256'h7D8A96959494929292939494919397847D95988684A38B8A7E869A9193929293),
    .INIT_69(256'h94928E9098837B95949297979494949595949493929292929192929393939796),
    .INIT_6A(256'h958F93929394969282899294938F9290988B8080808080808080808080939D98),
    .INIT_6B(256'h9190908F909091929591987F7C989593868C84898D7F9F959492929393949393),
    .INIT_6C(256'h938080829492948E91929393939393939392929292929292938D939892909393),
    .INIT_6D(256'h93929482869491959087938E9589808080808080808080808088979895959391),
    .INIT_6E(256'h8F909092969398837E9492988F7B8EA19C828194939292939393939392919292),
    .INIT_6F(256'h968D909090919192929292929191919292939393928E92909392949290908F8E),
    .INIT_70(256'h829690948980969297898080808080808080808080808596959593939798848D),
    .INIT_71(256'h91979383859495978777859D9684829292919293939292928F9291929391927D),
    .INIT_72(256'h90919191919190908F8F9092939395949191948F969495919190909090919192),
    .INIT_73(256'h85819996968D8080808080808080808080808295908F91919092837E9399928E),
    .INIT_74(256'h929496958D8898919E827D979291929293929292929392919391937D80979094),
    .INIT_75(256'h9191919191919191929394949390939396939492929191919192929292948386),
    .INIT_76(256'h92958980808080808080808080808C958C8E929191989C8383908D9291919191),
    .INIT_77(256'h82849A90927F86929392929393939393939192909292927F819A939586849794),
    .INIT_78(256'h94939292919191929490939392929594939292929293939495937D8894919296),
    .INIT_79(256'h808080808080808080808F978E8F93959494977E839796919292929394949595),
    .INIT_7A(256'h92938287969494959595959495919593959693808399949685859591919B9380),
    .INIT_7B(256'h949493959597999795999B96989797979798989894998B869192939487809797),
    .INIT_7C(256'h808080808080879893929096969498818495988E929293949596969797969595),
    .INIT_7D(256'h9A9797989898989797949797969A97827C97977E7C809998949A938080808080),
    .INIT_7E(256'h8B8C8C8C8D8D8D8D8C8C8C8C8C8D8E8A9A978D9092959194828396909498878B),
    .INIT_7F(256'h8080869C9A929297919695978A819893949294969694949897969B9C80858C8B),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_5000x8_sub_000000_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(addra[12]),
    .dia({open_n51,open_n52,open_n53,open_n54,open_n55,open_n56,open_n57,open_n58,8'b00000000}),
    .rsta(rsta),
    .doa({open_n80,open_n81,open_n82,open_n83,open_n84,open_n85,open_n86,open_n87,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=4096;data_offset=0;depth=904;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=4096;working_width=8;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h888989888A8A8A868B9FA0878E9A978C80A0A2969A9988808080808080808080),
    .INIT_01(256'h808080808080808080808080878A8090899B989D8E8A9A95919B96808B888888),
    .INIT_02(256'h979996959496909A878A9B9696989486808689878B898A8A8080808080808080),
    .INIT_03(256'h80808080809096808093978F808D8C87989EA19580808080808080808080808A),
    .INIT_04(256'h8080808080808080808080808090898B808F9C9E8B9580808080808080808080),
    .INIT_05(256'h989295A096929D8A8F958B808080808080808080808080808080808080808080),
    .INIT_06(256'h8080808080808080808080808A8D9080808080808080808080808080909B9793),
    .INIT_07(256'h80808080808080808080808080808E8E80808080808080808080808080808080),
    .INIT_08(256'h8095888280808080808080808080808080808080808080808080808080808080),
    .INIT_09(256'h808080808080808080808080808080808080808080808080878F8B8685858E80),
    .INIT_0A(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0C(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0D(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0E(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_0F(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_10(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_11(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_12(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_13(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_14(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_15(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_16(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_17(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_18(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_19(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1A(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1B(256'h8080808080808080808080808080808080808080808080808080808080808080),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000008080808080808080),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_5000x8_sub_004096_000 (
    .addra(addra[11:1]),
    .addrb(11'b00000000000),
    .bytea(addra[0]),
    .byteb(1'b0),
    .clka(clka),
    .csa(addra[12]),
    .dia({open_n108,open_n109,open_n110,open_n111,open_n112,open_n113,open_n114,open_n115,8'b00000000}),
    .rsta(rsta),
    .doa({open_n137,open_n138,open_n139,open_n140,open_n141,open_n142,open_n143,open_n144,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped),
    .o(doa[7]));

endmodule 

